netcdf SpringNetwork {

dimensions:
	spatialdim = 3;
	particle_number = 174;
	particlename_length = 5;
	chainname_length = 4;
	resname_length = 4;

	springdim = 2; 
	spring_number = 993;

variables:
	float   coordinates(particle_number, spatialdim); 
	        coordinates:units = "angstrom" ;
	        coordinates:long_name = "Particle coordinates";

	int     particleids(particle_number); 
	        particleids:long_name = "Particle ids in source database";

	char    particlenames(particle_number,particlename_length); 
	        particlenames:long_name = "Particle name";

	float   charges(particle_number);
	        charges:long_name = "Particle charge id";
	        charges:units = "electron" ;

	float   radii(particle_number);
	        radii:units = "A" ;
	        radii:long_name = "Particle radius";

	float   epsilon(particle_number);
	        epsilon:units = "kJ.mol-1" ;
	        epsilon:long_name = "Particle epsilon for Lennard-Jones";

	float   mass(particle_number);
	        mass:units = "Da" ;
	        mass:long_name = "Particle mass";

	float   surfaceaccessibility(particle_number);
	        surfaceaccessibility:units = "A2 or percent" ;
	        surfaceaccessibility:long_name = "Particle surface accessibility";

	float   hydrophobicityscale(particle_number);
	        hydrophobicityscale:units = "kJ.mol-1" ;
	        hydrophobicityscale:long_name = "Particle hydrophobicity scale (transfer energy)";

	char    resnames(particle_number,resname_length); 
	        resnames:long_name = "particle residue name";

	int     resids(particle_number); 
	        resids:long_name = "particle residue id";

	char    chainnames(particle_number,chainname_length); 
	        chainnames:long_name = "Chain name ";

	byte    dynamicstate(particle_number); 
	        dynamicstate:long_name = "particle dynamic state (static 0 or dynamic 1)";

	int     nbspringsperparticle(particle_number); 
	        nbspringsperparticle:long_name = "Number of springs per particle";

	int     springs(spring_number,springdim); 
	        springs:long_name = "Spring between particle referenced by 2 particle ids"; 

	float   springsstiffness(spring_number); 
	        springsstiffness:long_name = "Spring stiffness";
	float   springsequilibrium(spring_number); 
	        springsequilibrium:long_name = "Spring distance equilibrium";
data:
	particleids = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	coordinates = 
9.27257, 34.0063, 15.0073,
10.826, 29.9497, 14.937,
14.3379, 32.3195, 12.3651,
16.3871, 27.5676, 14.4209,
19.985, 30.2409, 15.4413,
22.8017, 26.984, 14.4686,
25.7259, 30.35, 16.929,
32.6787, 29.158, 14.972,
35.7699, 30.3063, 15.2976,
37.6656, 32.2484, 20.7806,
34.8493, 34.0841, 18.1909,
32.578, 34.8545, 21.299,
30.101, 30.8927, 20.5457,
29.6876, 36.4533, 24.94,
26.8071, 36.4533, 21.56,
24.7861, 32.9681, 23.414,
25.5082, 35.9865, 28.7448,
23.2475, 38.6895, 24.775,
20.9878, 36.4891, 22.1399,
19.7917, 32.6722, 27.1954,
20.6584, 38.6414, 28.7202,
19.4335, 41.9021, 24.6698,
15.2835, 37.0991, 23.416,
13.2723, 36.6217, 27.4599,
10.8033, 33.7516, 24.4406,
15.2975, 32.2915, 23.3545,
14.6393, 26.7528, 23.1978,
19.9474, 27.5401, 24.843,
19.8884, 22.7739, 27.0603,
21.987, 16.196, 26.5436,
24.3407, 14.5151, 29.4147,
25.497, 10.518, 29.6977,
27.4255, 14.8075, 33.3431,
26.226, 12.9474, 36.4524,
24.725, 15.4484, 38.2364,
29.1182, 19.298, 37.3449,
27.4427, 19.4937, 42.8023,
23.5243, 21.784, 41.8913,
24.2172, 20.6993, 37.8339,
19.1669, 21.8646, 37.5831,
17.2479, 18.3076, 34.7534,
17.4062, 21.3493, 31.9398,
18.6823, 24.3683, 33.583,
22.5823, 23.057, 33.7578,
24.0567, 19.7922, 30.4262,
18.1955, 17.8503, 29.2456,
21.4328, 15.6383, 33.749,
19.7389, 11.1943, 29.8776,
20.6864, 6.34675, 30.8195,
23.5844, 5.986, 28.9946,
20.8526, 3.17443, 27.0321,
16.2348, 7.46782, 26.2682,
22.1576, 9.95064, 24.3092,
22.291, 4.88578, 21.5724,
17.3317, 4.114, 22.9983,
17.1339, 9.19938, 21.6706,
21.2996, 8.24675, 18.5569,
19.1558, 4.5695, 17.1185,
14.5572, 6.86144, 18.0778,
16.4615, 10.7615, 15.6343,
14.6976, 12.0587, 18.5444,
19.934, 13.3175, 18.9741,
19.4709, 17.3528, 15.8631,
24.2418, 17.1602, 17.7352,
26.5438, 11.739, 18.8669,
29.2836, 13.9096, 21.0648,
31.7813, 10.6176, 22.3879,
32.4225, 14.2346, 25.783,
35.909, 14.4347, 28.665,
36.9147, 10.1093, 25.2603,
33.9762, 8.676, 26.078,
33.9318, 9.47462, 30.2506,
30.5587, 12.3059, 28.9038,
27.7259, 9.50909, 24.361,
23.447, 16.6658, 22.833,
21.0453, 18.6999, 20.3523,
17.4164, 16.777, 22.4726,
14.7554, 17.3402, 18.7554,
11.6397, 16.0254, 21.4696,
13.083, 20.4594, 22.5664,
13.899, 22.3554, 18.7237,
10.9535, 20.2382, 15.1923,
8.2396, 22.4366, 20.148,
9.5892, 25.6502, 19.7682,
9.0538, 25.8148, 16.2822,
5.6428, 24.7654, 16.6436,
5.06357, 27.0519, 19.6491,
6.85775, 30.1823, 17.7302,
9.18143, 30.0831, 20.2727,
12.5033, 31.8569, 19.4676,
15.549, 28.4306, 18.7414,
20.0191, 29.782, 20.4755,
21.3995, 25.7996, 18.843,
26.3921, 27.0797, 21.7803,
27.2724, 24.0217, 18.1213,
30.9526, 22.227, 16.4964,
31.7725, 23.9569, 12.6406,
30.0242, 19.51, 13.176,
27.0128, 20.1833, 14.5343,
26.0454, 22.549, 12.565,
28.0243, 20.2261, 8.15764,
24.2486, 17.8532, 11.6352,
21.655, 20.5879, 13.2451,
21.1074, 22.2953, 7.77422,
22.4226, 16.6264, 7.394,
18.3236, 16.7671, 11.1887,
15.9396, 21.2014, 11.4085,
16.7347, 21.4827, 6.95671,
13.8909, 23.772, 8.85944,
17.7322, 25.7674, 10.1356,
19.7729, 29.259, 10.2657,
23.8683, 27.9254, 9.84943,
25.1039, 31.6296, 12.2817,
30.915, 31.6185, 10.9344,
30.573, 34.5413, 15.1699,
33.402, 36.3244, 12.8036,
36.6611, 37.3569, 13.4354,
37.4493, 41.2741, 13.8906,
44.1064, 35.1571, 11.8332,
46.2171, 40.6596, 13.5792,
42.0645, 40.0154, 17.1658,
41.5218, 35.2044, 16.6691,
46.9572, 35.4206, 15.5557,
46.434, 37.5302, 19.5506,
41.9072, 36.9629, 21.0205,
44.5199, 32.1247, 20.1539,
49.1802, 34.06, 21.2559,
48.266, 35.6332, 24.5585,
49.5555, 37.9561, 28.3077,
52.6345, 33.1087, 26.0245,
51.95, 31.2531, 28.9109,
50.2699, 27.7196, 25.6978,
53.8353, 25.7527, 24.4676,
54.4046, 27.35, 20.6594,
53.2772, 23.0706, 19.7156,
49.8296, 24.245, 21.6901,
49.9959, 28.6246, 20.3859,
51.0624, 27.0277, 15.5391,
46.5178, 21.7872, 18.1956,
44.9608, 26.7786, 20.4908,
46.9474, 29.5276, 15.096,
45.9125, 24.8289, 12.1709,
42.3983, 24.7829, 14.3124,
41.5082, 28.6544, 13.2942,
44.2276, 30.3499, 8.71455,
40.6845, 24.6595, 9.6415,
37.553, 26.8542, 12.9288,
38.0903, 30.9819, 9.60213,
36.9848, 27.9116, 5.9996,
33.395, 27.2694, 6.9644,
33.0622, 31.8202, 6.33556,
30.5993, 29.5665, 3.06375,
28.7676, 25.803, 4.09825,
27.8394, 28.261, 8.14382,
23.0222, 29.6459, 6.067,
23.2497, 34.0417, 7.33022,
28.1223, 35.6089, 8.39,
27.9454, 37.7721, 12.2477,
31.4313, 40.4811, 12.0044,
32.3047, 39.8986, 17.0999,
33.4888, 44.3316, 13.4081,
31.1475, 46.3913, 20.737,
29.1469, 41.7795, 22.1991,
27.2734, 45.129, 22.5544,
26.4636, 41.2746, 17.0808,
23.6752, 40.6985, 19.6947,
21.6726, 43.0094, 17.5042,
23.4756, 41.5076, 13.1856,
21.9166, 37.374, 15.8504,
17.976, 40.0223, 17.6967,
18.0501, 36.2669, 12.3044,
16.2684, 35.1711, 16.4154,
12.8297, 38.3559, 16.5859,
13.6722, 41.3877, 13.838;
	charges = 
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
1,
0,
0,
1,
-1,
1,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
1,
0,
0,
1,
0,
0,
-1,
0,
-1,
0,
0,
-1,
0,
1,
0,
0,
-1,
0,
0,
1,
0,
0,
0,
0,
0,
-1,
0,
0,
-1,
0,
0,
-1,
0,
0,
-1,
0,
1,
0,
0,
0,
1,
1,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
-1,
0,
0,
0,
0,
1,
0,
0,
1,
1,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
1,
0,
0,
0,
1,
0,
0,
-1,
0,
0,
-1,
0,
0,
0,
1,
1,
0,
-1,
0,
0,
1,
0,
-1,
0,
0,
0,
0,
0,
-1,
0,
-1,
1,
0,
0,
0,
0,
1,
1,
0,
-1,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0;
	radii = 
3.3,
2.58,
3.47,
3.3,
3.3,
3.3,
3.49,
2.58,
3.2,
2.88,
3.3,
2.58,
3.44,
3.12,
3.3,
3.3,
3.47,
3.03,
3.49,
3.47,
3.22,
3.47,
3.47,
3.2,
3.13,
3.49,
3.38,
3.64,
3.3,
2.88,
3.12,
3.12,
3.47,
2.88,
3.2,
3.47,
3.2,
2.58,
3.22,
3.3,
3,
2.58,
3.3,
3,
3.66,
3.38,
3.64,
3.47,
3,
3.2,
3.12,
3.47,
3.64,
3.34,
3.34,
3.49,
3.47,
3,
3.34,
2.58,
3.22,
3.49,
3.49,
3.22,
3.85,
2.88,
3.22,
3.47,
3.38,
2.58,
2.58,
3.49,
3.38,
3.47,
2.58,
3.12,
3.49,
2.88,
3.34,
3.2,
3.3,
3.47,
2.88,
2.88,
2.88,
2.88,
3.12,
2.58,
3.3,
3.2,
3.3,
3.49,
3.47,
3.22,
3.3,
3,
3.49,
2.88,
2.58,
2.88,
3.47,
2.88,
3.47,
3.44,
3.44,
3.12,
3.47,
3.2,
3.22,
2.88,
3.3,
3.12,
3.3,
3.64,
3.49,
2.88,
3.2,
3.2,
3.85,
3.34,
3,
3.49,
3.34,
2.88,
3.47,
3.49,
3.47,
2.58,
3.47,
2.58,
3.12,
3.22,
3.12,
2.88,
3,
3.3,
3.47,
3.34,
3.47,
3.47,
3.49,
3,
3.12,
2.88,
3.47,
3.47,
3.22,
3.49,
2.88,
2.88,
3.34,
2.58,
3,
3.64,
3,
3.44,
3.3,
3.3,
3.3,
3.13,
3.47,
3.47,
3.49,
3.22,
2.88,
3.03,
2.88,
3.22,
3.49,
3.3,
3.49,
3.49,
3.3,
2.58;
	epsilon = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	mass = 
117,
75,
174,
117,
117,
117,
131,
75,
115,
89,
117,
75,
146,
119,
117,
117,
174,
121,
131,
174,
147,
174,
131,
115,
132,
131,
155,
165,
117,
89,
119,
119,
174,
89,
115,
174,
115,
75,
147,
117,
133,
75,
117,
133,
181,
155,
165,
131,
133,
115,
119,
174,
165,
146,
146,
131,
131,
133,
146,
75,
147,
131,
131,
147,
204,
89,
147,
131,
155,
75,
75,
131,
155,
174,
75,
119,
131,
89,
146,
115,
117,
174,
89,
89,
89,
89,
119,
75,
117,
115,
117,
131,
131,
147,
117,
133,
131,
89,
75,
89,
174,
89,
131,
146,
146,
119,
149,
115,
147,
89,
117,
119,
117,
165,
131,
89,
115,
115,
204,
146,
133,
131,
146,
89,
174,
131,
131,
75,
174,
75,
119,
147,
119,
89,
133,
117,
131,
146,
174,
174,
131,
133,
119,
89,
174,
131,
147,
131,
89,
89,
146,
75,
133,
165,
133,
146,
117,
117,
117,
132,
174,
174,
131,
147,
89,
121,
89,
147,
131,
117,
131,
131,
117,
75;
	surfaceaccessibility = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	hydrophobicityscale = 
5.04836,
0,
-4.17938,
5.04836,
5.04836,
5.04836,
7.0346,
0,
2.97936,
1.28278,
5.04836,
0,
-4.09662,
1.07588,
5.04836,
5.04836,
-4.17938,
6.37252,
7.0346,
-4.17938,
-2.64832,
-4.17938,
7.4484,
2.97936,
-2.4828,
7.0346,
0.53794,
7.40702,
5.04836,
1.28278,
1.07588,
1.07588,
-4.17938,
1.28278,
2.97936,
-4.17938,
2.97936,
0,
-2.64832,
5.04836,
-3.18626,
0,
5.04836,
-3.18626,
3.97248,
0.53794,
7.40702,
7.4484,
-3.18626,
2.97936,
1.07588,
-4.17938,
7.40702,
-0.91036,
-0.91036,
7.0346,
7.4484,
-3.18626,
-0.91036,
0,
-2.64832,
7.0346,
7.0346,
-2.64832,
9.3105,
1.28278,
-2.64832,
7.4484,
0.53794,
0,
0,
7.0346,
0.53794,
-4.17938,
0,
1.07588,
7.0346,
1.28278,
-0.91036,
2.97936,
5.04836,
-4.17938,
1.28278,
1.28278,
1.28278,
1.28278,
1.07588,
0,
5.04836,
2.97936,
5.04836,
7.0346,
7.4484,
-2.64832,
5.04836,
-3.18626,
7.0346,
1.28278,
0,
1.28278,
-4.17938,
1.28278,
7.4484,
-4.09662,
-4.09662,
1.07588,
5.08974,
2.97936,
-2.64832,
1.28278,
5.04836,
1.07588,
5.04836,
7.40702,
7.0346,
1.28278,
2.97936,
2.97936,
9.3105,
-0.91036,
-3.18626,
7.0346,
-0.91036,
1.28278,
-4.17938,
7.0346,
7.4484,
0,
-4.17938,
0,
1.07588,
-2.64832,
1.07588,
1.28278,
-3.18626,
5.04836,
7.4484,
-0.91036,
-4.17938,
-4.17938,
7.0346,
-3.18626,
1.07588,
1.28278,
-4.17938,
7.4484,
-2.64832,
7.0346,
1.28278,
1.28278,
-0.91036,
0,
-3.18626,
7.40702,
-3.18626,
-4.09662,
5.04836,
5.04836,
5.04836,
-2.4828,
-4.17938,
-4.17938,
7.0346,
-2.64832,
1.28278,
6.37252,
1.28278,
-2.64832,
7.0346,
5.04836,
7.0346,
7.0346,
5.04836,
0;
	particlenames = 
"VCA",
"GCA",
"RCA",
"VCA",
"VCA",
"VCA",
"LCA",
"GCA",
"PCA",
"ACA",
"VCA",
"GCA",
"KCA",
"TCA",
"VCA",
"VCA",
"RCA",
"CCA",
"LCA",
"RCA",
"ECA",
"RCA",
"ICA",
"PCA",
"NCA",
"LCA",
"HCA",
"FCA",
"VCA",
"ACA",
"TCA",
"TCA",
"RCA",
"ACA",
"PCA",
"RCA",
"PCA",
"GCA",
"ECA",
"VCA",
"DCA",
"GCA",
"VCA",
"DCA",
"YCA",
"HCA",
"FCA",
"ICA",
"DCA",
"PCA",
"TCA",
"RCA",
"FCA",
"QCA",
"QCA",
"LCA",
"ICA",
"DCA",
"QCA",
"GCA",
"ECA",
"LCA",
"LCA",
"ECA",
"WCA",
"ACA",
"ECA",
"ICA",
"HCA",
"GCA",
"GCA",
"LCA",
"HCA",
"RCA",
"GCA",
"TCA",
"LCA",
"ACA",
"QCA",
"PCA",
"VCA",
"RCA",
"ACA",
"ACA",
"ACA",
"ACA",
"TCA",
"GCA",
"VCA",
"PCA",
"VCA",
"LCA",
"ICA",
"ECA",
"VCA",
"DCA",
"LCA",
"ACA",
"GCA",
"ACA",
"RCA",
"ACA",
"ICA",
"KCA",
"KCA",
"TCA",
"MCA",
"PCA",
"ECA",
"ACA",
"VCA",
"TCA",
"VCA",
"FCA",
"LCA",
"ACA",
"PCA",
"PCA",
"WCA",
"QCA",
"DCA",
"LCA",
"QCA",
"ACA",
"RCA",
"LCA",
"ICA",
"GCA",
"RCA",
"GCA",
"TCA",
"ECA",
"TCA",
"ACA",
"DCA",
"VCA",
"ICA",
"QCA",
"RCA",
"RCA",
"LCA",
"DCA",
"TCA",
"ACA",
"RCA",
"ICA",
"ECA",
"LCA",
"ACA",
"ACA",
"QCA",
"GCA",
"DCA",
"FCA",
"DCA",
"KCA",
"VCA",
"VCA",
"VCA",
"NCA",
"RCA",
"RCA",
"LCA",
"ECA",
"ACA",
"CCA",
"ACA",
"ECA",
"LCA",
"VCA",
"LCA",
"LCA",
"VCA",
"GCA";
	resnames = 
"VAL",
"GLY",
"ARG",
"VAL",
"VAL",
"VAL",
"LEU",
"GLY",
"PRO",
"ALA",
"VAL",
"GLY",
"LYS",
"THR",
"VAL",
"VAL",
"ARG",
"CYS",
"LEU",
"ARG",
"GLU",
"ARG",
"ILE",
"PRO",
"ASN",
"LEU",
"HIS",
"PHE",
"VAL",
"ALA",
"THR",
"THR",
"ARG",
"ALA",
"PRO",
"ARG",
"PRO",
"GLY",
"GLU",
"VAL",
"ASP",
"GLY",
"VAL",
"ASP",
"TYR",
"HIS",
"PHE",
"ILE",
"ASP",
"PRO",
"THR",
"ARG",
"PHE",
"GLN",
"GLN",
"LEU",
"ILE",
"ASP",
"GLN",
"GLY",
"GLU",
"LEU",
"LEU",
"GLU",
"TRP",
"ALA",
"GLU",
"ILE",
"HIS",
"GLY",
"GLY",
"LEU",
"HIS",
"ARG",
"GLY",
"THR",
"LEU",
"ALA",
"GLN",
"PRO",
"VAL",
"ARG",
"ALA",
"ALA",
"ALA",
"ALA",
"THR",
"GLY",
"VAL",
"PRO",
"VAL",
"LEU",
"ILE",
"GLU",
"VAL",
"ASP",
"LEU",
"ALA",
"GLY",
"ALA",
"ARG",
"ALA",
"ILE",
"LYS",
"LYS",
"THR",
"MET",
"PRO",
"GLU",
"ALA",
"VAL",
"THR",
"VAL",
"PHE",
"LEU",
"ALA",
"PRO",
"PRO",
"TRP",
"GLN",
"ASP",
"LEU",
"GLN",
"ALA",
"ARG",
"LEU",
"ILE",
"GLY",
"ARG",
"GLY",
"THR",
"GLU",
"THR",
"ALA",
"ASP",
"VAL",
"ILE",
"GLN",
"ARG",
"ARG",
"LEU",
"ASP",
"THR",
"ALA",
"ARG",
"ILE",
"GLU",
"LEU",
"ALA",
"ALA",
"GLN",
"GLY",
"ASP",
"PHE",
"ASP",
"LYS",
"VAL",
"VAL",
"VAL",
"ASN",
"ARG",
"ARG",
"LEU",
"GLU",
"ALA",
"CYS",
"ALA",
"GLU",
"LEU",
"VAL",
"LEU",
"LEU",
"VAL",
"GLY";
	resids = 
1,
2,
3,
4,
5,
6,
7,
9,
10,
12,
13,
14,
15,
17,
18,
19,
20,
21,
22,
23,
24,
25,
26,
27,
28,
29,
30,
31,
33,
35,
36,
37,
38,
39,
40,
41,
42,
43,
44,
45,
46,
47,
48,
49,
50,
51,
52,
53,
54,
55,
56,
57,
58,
59,
60,
61,
62,
63,
64,
65,
66,
67,
68,
69,
70,
71,
72,
73,
74,
75,
76,
77,
78,
79,
81,
82,
83,
84,
85,
86,
87,
88,
89,
90,
91,
92,
93,
94,
95,
96,
97,
98,
99,
100,
101,
102,
103,
104,
105,
106,
107,
108,
109,
110,
111,
112,
113,
114,
115,
116,
117,
118,
119,
120,
121,
122,
123,
124,
126,
127,
128,
129,
130,
131,
132,
133,
134,
135,
136,
137,
138,
139,
140,
141,
142,
143,
144,
145,
146,
147,
148,
149,
150,
151,
152,
153,
154,
155,
156,
157,
158,
159,
160,
161,
162,
163,
164,
165,
166,
167,
168,
169,
170,
171,
173,
174,
175,
176,
177,
178,
180,
181,
182,
183;
	chainnames = 
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"",
"";
	dynamicstate = 
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1;
	nbspringsperparticle = 
9,
13,
11,
19,
15,
18,
16,
17,
15,
8,
14,
12,
12,
9,
15,
14,
7,
15,
16,
11,
8,
9,
12,
6,
7,
12,
16,
9,
13,
14,
15,
13,
11,
8,
11,
8,
4,
6,
12,
9,
10,
9,
8,
11,
15,
13,
14,
12,
7,
10,
8,
9,
18,
11,
10,
15,
11,
8,
9,
9,
10,
16,
15,
15,
10,
9,
9,
10,
6,
6,
8,
9,
12,
14,
14,
15,
15,
14,
8,
11,
16,
10,
12,
14,
14,
9,
8,
11,
13,
18,
17,
15,
15,
9,
14,
9,
12,
9,
12,
16,
12,
11,
19,
14,
9,
12,
14,
8,
8,
12,
15,
17,
15,
21,
16,
15,
14,
9,
11,
6,
9,
15,
12,
9,
9,
13,
13,
9,
4,
8,
6,
10,
7,
8,
7,
9,
14,
8,
8,
11,
14,
9,
10,
14,
10,
8,
13,
15,
10,
12,
9,
8,
8,
16,
11,
9,
13,
13,
11,
14,
8,
5,
10,
8,
16,
12,
11,
9,
13,
13,
11,
16,
9,
6;
	springs = 
0, 1,
0, 84,
0, 88,
0, 87,
0, 89,
0, 172,
0, 173,
0, 2,
0, 171,
1, 83,
1, 84,
1, 85,
1, 86,
1, 88,
1, 87,
1, 89,
1, 172,
1, 3,
1, 90,
1, 2,
1, 171,
2, 89,
2, 172,
2, 109,
2, 110,
2, 3,
2, 90,
2, 4,
2, 170,
2, 171,
3, 108,
3, 80,
3, 83,
3, 84,
3, 89,
3, 102,
3, 106,
3, 109,
3, 110,
3, 5,
3, 90,
3, 91,
3, 92,
3, 26,
3, 4,
3, 171,
3, 111,
4, 89,
4, 109,
4, 110,
4, 5,
4, 90,
4, 91,
4, 92,
4, 168,
4, 170,
4, 171,
4, 111,
4, 6,
4, 112,
5, 102,
5, 103,
5, 109,
5, 110,
5, 154,
5, 90,
5, 91,
5, 92,
5, 98,
5, 111,
5, 153,
5, 94,
5, 99,
5, 93,
5, 6,
5, 112,
6, 91,
6, 92,
6, 168,
6, 111,
6, 94,
6, 99,
6, 93,
6, 113,
6, 12,
6, 112,
6, 114,
6, 14,
6, 15,
6, 7,
7, 153,
7, 94,
7, 95,
7, 96,
7, 113,
7, 12,
7, 112,
7, 114,
7, 149,
7, 146,
7, 147,
7, 8,
7, 9,
7, 10,
7, 115,
7, 11,
8, 96,
8, 113,
8, 12,
8, 114,
8, 146,
8, 147,
8, 9,
8, 10,
8, 115,
8, 116,
8, 11,
8, 142,
8, 143,
8, 121,
9, 12,
9, 10,
9, 11,
9, 121,
9, 124,
9, 125,
10, 113,
10, 12,
10, 114,
10, 13,
10, 115,
10, 116,
10, 11,
10, 117,
10, 159,
10, 121,
10, 124,
11, 12,
11, 114,
11, 13,
11, 14,
11, 15,
11, 162,
11, 115,
11, 159,
12, 94,
12, 93,
12, 114,
12, 13,
12, 14,
12, 15,
13, 14,
13, 15,
13, 16,
13, 17,
13, 162,
13, 159,
14, 168,
14, 18,
14, 114,
14, 15,
14, 16,
14, 17,
14, 164,
14, 165,
14, 162,
14, 163,
14, 159,
15, 91,
15, 27,
15, 18,
15, 19,
15, 20,
15, 93,
15, 16,
15, 17,
15, 165,
16, 18,
16, 19,
16, 20,
16, 17,
17, 18,
17, 19,
17, 20,
17, 22,
17, 166,
17, 169,
17, 21,
17, 164,
17, 165,
17, 162,
17, 163,
18, 91,
18, 168,
18, 171,
18, 19,
18, 20,
18, 22,
18, 25,
18, 166,
18, 169,
18, 21,
18, 164,
18, 165,
19, 23,
19, 91,
19, 26,
19, 27,
19, 20,
19, 22,
19, 25,
20, 23,
20, 22,
20, 21,
21, 23,
21, 22,
21, 166,
21, 169,
21, 165,
21, 163,
22, 89,
22, 172,
22, 23,
22, 24,
22, 171,
22, 25,
22, 169,
23, 24,
23, 25,
24, 88,
24, 87,
24, 89,
24, 26,
24, 25,
25, 88,
25, 89,
25, 90,
25, 91,
25, 26,
25, 27,
25, 171,
26, 79,
26, 80,
26, 82,
26, 83,
26, 84,
26, 88,
26, 89,
26, 90,
26, 91,
26, 92,
26, 27,
26, 28,
27, 90,
27, 91,
27, 92,
27, 28,
27, 93,
28, 79,
28, 75,
28, 29,
28, 45,
28, 76,
28, 92,
28, 41,
28, 42,
28, 43,
28, 74,
28, 44,
29, 47,
29, 52,
29, 61,
29, 75,
29, 45,
29, 76,
29, 46,
29, 41,
29, 31,
29, 30,
29, 74,
29, 32,
29, 44,
30, 47,
30, 52,
30, 45,
30, 46,
30, 31,
30, 49,
30, 73,
30, 72,
30, 74,
30, 32,
30, 33,
30, 34,
30, 44,
30, 67,
31, 47,
31, 52,
31, 48,
31, 46,
31, 49,
31, 73,
31, 72,
31, 32,
31, 33,
31, 71,
31, 67,
32, 46,
32, 72,
32, 33,
32, 34,
32, 35,
32, 38,
32, 44,
32, 71,
33, 46,
33, 72,
33, 34,
33, 35,
33, 38,
34, 40,
34, 46,
34, 39,
34, 35,
34, 38,
34, 44,
34, 36,
34, 37,
35, 43,
35, 38,
35, 44,
35, 36,
35, 37,
36, 38,
36, 37,
37, 39,
37, 43,
37, 38,
38, 40,
38, 46,
38, 39,
38, 42,
38, 43,
38, 44,
39, 40,
39, 46,
39, 41,
39, 42,
39, 43,
39, 44,
40, 47,
40, 45,
40, 46,
40, 41,
40, 42,
40, 43,
40, 44,
41, 45,
41, 46,
41, 42,
41, 43,
41, 44,
42, 45,
42, 43,
42, 44,
43, 45,
43, 46,
43, 44,
44, 45,
44, 46,
44, 74,
45, 79,
45, 47,
45, 76,
45, 46,
45, 74,
46, 47,
47, 50,
47, 51,
47, 52,
47, 55,
47, 48,
47, 49,
48, 50,
48, 51,
48, 52,
48, 54,
48, 49,
49, 50,
49, 51,
49, 52,
49, 53,
49, 54,
49, 73,
50, 51,
50, 52,
50, 53,
50, 54,
50, 55,
51, 58,
51, 52,
51, 53,
51, 54,
51, 55,
52, 56,
52, 53,
52, 54,
52, 55,
52, 61,
52, 76,
52, 64,
52, 73,
52, 65,
52, 74,
53, 56,
53, 57,
53, 58,
53, 54,
53, 55,
53, 64,
53, 73,
54, 56,
54, 57,
54, 58,
54, 55,
55, 78,
55, 56,
55, 57,
55, 58,
55, 59,
55, 60,
55, 61,
55, 77,
55, 76,
56, 57,
56, 58,
56, 59,
56, 60,
56, 61,
56, 64,
56, 73,
57, 58,
57, 59,
57, 60,
57, 61,
58, 59,
58, 60,
58, 61,
59, 60,
59, 105,
59, 61,
59, 62,
59, 77,
60, 78,
60, 61,
60, 62,
60, 77,
60, 76,
61, 105,
61, 62,
61, 75,
61, 77,
61, 76,
61, 64,
61, 63,
61, 74,
62, 80,
62, 104,
62, 105,
62, 75,
62, 77,
62, 102,
62, 76,
62, 106,
62, 101,
62, 63,
62, 98,
62, 74,
63, 105,
63, 75,
63, 102,
63, 76,
63, 64,
63, 101,
63, 97,
63, 98,
63, 65,
63, 74,
63, 94,
63, 95,
63, 99,
64, 75,
64, 66,
64, 73,
64, 65,
64, 74,
65, 66,
65, 73,
65, 72,
65, 74,
65, 70,
65, 67,
66, 73,
66, 72,
66, 69,
66, 70,
66, 71,
66, 67,
66, 68,
67, 73,
67, 72,
67, 69,
67, 70,
67, 71,
67, 68,
68, 72,
68, 69,
68, 70,
68, 71,
69, 72,
69, 70,
69, 71,
70, 73,
70, 72,
70, 71,
71, 73,
71, 72,
72, 73,
73, 74,
74, 75,
74, 76,
75, 79,
75, 80,
75, 77,
75, 102,
75, 76,
75, 92,
75, 98,
75, 94,
76, 78,
76, 79,
76, 80,
76, 77,
77, 81,
77, 78,
77, 79,
77, 80,
77, 82,
77, 105,
77, 106,
78, 81,
78, 79,
78, 80,
78, 82,
79, 81,
79, 80,
79, 82,
79, 83,
80, 81,
80, 82,
80, 83,
80, 84,
80, 85,
80, 106,
80, 90,
80, 92,
81, 108,
81, 82,
81, 83,
81, 84,
81, 85,
81, 106,
82, 83,
82, 84,
82, 85,
82, 86,
82, 88,
82, 87,
83, 84,
83, 85,
83, 86,
83, 88,
83, 87,
83, 89,
83, 90,
84, 85,
84, 86,
84, 88,
84, 87,
84, 89,
84, 90,
85, 86,
85, 88,
85, 87,
86, 88,
86, 87,
86, 89,
87, 88,
87, 89,
87, 90,
88, 89,
88, 90,
89, 172,
89, 90,
89, 91,
89, 171,
90, 91,
90, 92,
90, 171,
91, 92,
91, 171,
91, 93,
92, 102,
92, 94,
92, 99,
92, 93,
93, 94,
93, 95,
94, 102,
94, 97,
94, 98,
94, 95,
94, 96,
94, 99,
95, 97,
95, 98,
95, 96,
95, 99,
95, 146,
96, 100,
96, 97,
96, 98,
96, 153,
96, 99,
96, 113,
96, 149,
96, 146,
97, 102,
97, 100,
97, 101,
97, 98,
97, 99,
98, 102,
98, 100,
98, 101,
98, 99,
99, 104,
99, 102,
99, 103,
99, 100,
99, 101,
99, 111,
99, 153,
100, 104,
100, 102,
100, 103,
100, 101,
100, 111,
100, 152,
100, 153,
100, 149,
101, 104,
101, 105,
101, 102,
101, 103,
101, 106,
102, 104,
102, 105,
102, 103,
102, 106,
102, 107,
102, 109,
102, 111,
103, 108,
103, 104,
103, 105,
103, 106,
103, 107,
103, 109,
103, 110,
103, 154,
103, 111,
104, 105,
104, 106,
104, 107,
105, 108,
105, 106,
105, 107,
106, 108,
106, 107,
106, 109,
106, 110,
107, 108,
107, 109,
107, 110,
108, 109,
108, 110,
109, 110,
109, 154,
109, 111,
110, 154,
110, 170,
110, 111,
110, 153,
110, 155,
110, 112,
111, 154,
111, 152,
111, 153,
111, 113,
111, 155,
111, 156,
111, 112,
112, 154,
112, 168,
112, 170,
112, 153,
112, 113,
112, 155,
112, 156,
112, 114,
112, 157,
113, 151,
113, 153,
113, 155,
113, 156,
113, 114,
113, 157,
113, 158,
113, 148,
113, 149,
113, 146,
113, 147,
113, 150,
113, 115,
113, 116,
114, 156,
114, 157,
114, 158,
114, 164,
114, 115,
114, 116,
114, 159,
115, 156,
115, 157,
115, 158,
115, 147,
115, 150,
115, 116,
115, 117,
115, 159,
115, 160,
116, 157,
116, 158,
116, 147,
116, 117,
116, 159,
116, 160,
116, 118,
116, 121,
116, 120,
117, 158,
117, 159,
117, 160,
117, 121,
117, 119,
117, 120,
118, 147,
118, 140,
118, 143,
118, 144,
118, 121,
118, 122,
118, 123,
118, 125,
118, 119,
118, 120,
119, 121,
119, 122,
119, 123,
119, 120,
120, 121,
120, 122,
120, 123,
120, 124,
120, 125,
121, 147,
121, 140,
121, 143,
121, 122,
121, 123,
121, 124,
121, 125,
122, 136,
122, 140,
122, 143,
122, 144,
122, 123,
122, 124,
122, 125,
122, 126,
123, 124,
123, 125,
123, 126,
123, 127,
124, 125,
124, 126,
124, 127,
125, 136,
125, 139,
125, 140,
125, 143,
125, 126,
125, 127,
126, 136,
126, 139,
126, 140,
126, 127,
126, 128,
126, 133,
126, 131,
126, 129,
126, 130,
127, 136,
127, 128,
127, 131,
127, 129,
127, 130,
128, 129,
128, 130,
129, 136,
129, 133,
129, 131,
129, 132,
129, 130,
130, 131,
130, 132,
131, 136,
131, 139,
131, 135,
131, 133,
131, 134,
131, 132,
132, 136,
132, 135,
132, 133,
132, 134,
133, 136,
133, 135,
133, 134,
133, 137,
134, 136,
134, 138,
134, 135,
134, 137,
135, 136,
135, 138,
135, 139,
135, 140,
135, 137,
136, 138,
136, 139,
136, 140,
136, 137,
137, 138,
137, 139,
137, 140,
137, 141,
138, 139,
138, 140,
138, 141,
138, 142,
139, 140,
139, 141,
139, 142,
139, 143,
140, 141,
140, 142,
140, 143,
140, 144,
141, 145,
141, 146,
141, 142,
141, 143,
141, 144,
142, 145,
142, 146,
142, 147,
142, 143,
142, 144,
143, 145,
143, 148,
143, 146,
143, 147,
143, 144,
144, 145,
144, 148,
144, 146,
144, 147,
145, 148,
145, 149,
145, 146,
145, 147,
146, 148,
146, 149,
146, 147,
147, 148,
147, 149,
147, 150,
148, 151,
148, 152,
148, 149,
148, 150,
149, 151,
149, 152,
149, 153,
149, 150,
150, 151,
150, 152,
150, 153,
150, 156,
151, 154,
151, 152,
151, 153,
151, 156,
152, 154,
152, 153,
153, 154,
153, 155,
153, 156,
154, 155,
154, 156,
155, 170,
155, 156,
155, 157,
156, 157,
156, 158,
156, 167,
157, 168,
157, 158,
157, 164,
157, 167,
157, 159,
157, 160,
158, 164,
158, 167,
158, 159,
158, 160,
159, 161,
159, 164,
159, 162,
159, 160,
160, 161,
160, 164,
161, 164,
161, 162,
161, 163,
162, 166,
162, 164,
162, 165,
162, 163,
163, 166,
163, 164,
163, 165,
164, 168,
164, 166,
164, 169,
164, 165,
164, 167,
165, 168,
165, 166,
165, 169,
165, 167,
166, 173,
166, 168,
166, 169,
166, 167,
167, 168,
167, 170,
167, 169,
168, 170,
168, 171,
168, 169,
169, 172,
169, 173,
169, 170,
169, 171,
170, 172,
170, 173,
170, 171,
171, 172,
171, 173,
172, 173;
	springsstiffness = 
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1;
	springsequilibrium = 
4.34437,
8.29299,
6.56689,
5.27912,
5.912,
5.83643,
8.67239,
5.95684,
7.23055,
6.58455,
4.69554,
7.52699,
7.98797,
5.585,
4.85832,
5.19388,
8.79751,
6.07186,
6.25206,
4.95622,
7.68556,
7.35018,
7.51842,
7.7086,
6.58126,
5.56837,
7.56628,
6.75822,
5.41901,
5.3163,
7.18101,
7.20221,
8.85903,
7.76625,
7.678,
8.8232,
7.05713,
4.83872,
5.62043,
6.44124,
4.48493,
7.39957,
6.9141,
8.9863,
4.59699,
7.86169,
8.7746,
8.64861,
7.29638,
5.27215,
4.41443,
5.81775,
5.0552,
5.77036,
7.40137,
7.06377,
6.25057,
7.19097,
5.93151,
6.17366,
6.61227,
8.34676,
6.77899,
5.65806,
8.81593,
8.54118,
7.18713,
4.7439,
7.99921,
4.83325,
8.18603,
6.48882,
5.81501,
8.14628,
5.09258,
5.62704,
6.74294,
6.56406,
8.0629,
7.71035,
6.62273,
8.9444,
5.88849,
8.02942,
5.70232,
4.86019,
6.64498,
7.73727,
7.05641,
7.32073,
8.41715,
8.09492,
7.30356,
5.77134,
5.0465,
6.38119,
8.40983,
5.78383,
8.25842,
5.76546,
7.83878,
3.31353,
8.25585,
6.27209,
7.52212,
8.51417,
7.95947,
6.658,
7.74741,
6.70511,
4.55055,
6.18698,
6.11794,
4.84673,
6.9314,
7.3466,
8.17871,
8.68417,
6.29848,
7.67833,
7.68872,
4.24363,
5.7397,
6.3649,
6.34627,
6.88398,
8.61481,
6.18683,
5.25565,
8.82083,
6.01132,
6.05042,
3.92591,
8.77203,
6.43996,
6.93487,
8.13067,
4.73277,
6.45634,
4.91605,
5.99392,
8.29124,
7.78065,
8.66091,
6.5689,
7.81591,
5.4607,
6.51415,
7.0994,
6.54208,
6.38613,
4.44086,
6.20475,
5.67113,
6.81926,
6.01442,
8.95475,
7.57395,
5.84832,
7.65972,
4.43486,
7.3162,
5.29225,
6.58987,
5.59559,
5.85247,
8.74496,
7.87317,
6.44288,
7.41078,
5.33371,
6.2714,
8.7966,
6.3184,
6.16845,
6.07895,
8.65021,
8.01949,
6.78702,
5.52893,
5.30812,
4.10999,
7.34906,
4.71914,
8.23417,
8.6027,
8.92565,
4.98779,
8.73079,
5.47985,
7.14044,
7.91241,
6.9781,
6.41901,
7.53522,
6.44651,
6.93123,
5.877,
7.17456,
8.02948,
6.42616,
6.17385,
8.85889,
5.56059,
7.62705,
7.31857,
8.80722,
5.64767,
6.22162,
7.36244,
5.92412,
7.76036,
7.70737,
5.34209,
8.58067,
6.4702,
7.58851,
7.36765,
6.64771,
8.73795,
7.12749,
7.36555,
4.54155,
5.68579,
7.32775,
4.80804,
6.96453,
4.84245,
6.30129,
5.78442,
8.56367,
5.58673,
8.07734,
4.8487,
7.19587,
4.80674,
6.02084,
6.07289,
5.57987,
6.81269,
7.57537,
6.51362,
6.31683,
8.29982,
6.20334,
8.93886,
7.03105,
6.67297,
4.84786,
6.74755,
8.09772,
5.61267,
7.63571,
7.57415,
4.90982,
6.41389,
5.25707,
7.15029,
8.47733,
7.93304,
6.92381,
5.64651,
7.94481,
8.88608,
5.65684,
6.82223,
7.22447,
8.23665,
6.13138,
6.41773,
6.63523,
8.35449,
6.74452,
4.94095,
6.14825,
7.24817,
8.75544,
7.38297,
4.07536,
4.01507,
8.81691,
5.68245,
5.69382,
7.18798,
6.99396,
5.33885,
4.17064,
8.57291,
7.87782,
6.61855,
6.9816,
5.00332,
7.45259,
8.87926,
5.38058,
8.86472,
5.80049,
6.36471,
6.46528,
7.69075,
4.96904,
5.87081,
5.42657,
5.95039,
7.21521,
8.517,
8.78071,
6.06356,
5.98183,
3.81658,
5.62566,
6.24859,
8.07306,
6.68614,
8.96294,
6.12566,
8.72727,
3.41919,
7.03501,
8.12626,
8.73007,
5.5688,
8.51391,
5.90881,
5.29074,
8.96186,
6.67813,
7.41209,
8.34962,
5.12076,
8.58674,
5.71213,
7.62506,
6.04502,
4.62923,
6.12806,
8.28624,
4.25663,
7.98634,
7.07485,
5.18911,
7.88459,
4.98464,
7.46479,
4.93375,
7.65519,
5.93407,
4.74389,
5.26502,
8.9122,
8.97653,
5.60738,
5.06438,
4.14645,
6.33711,
7.21134,
8.20294,
4.48598,
7.21816,
3.66648,
5.74565,
6.99596,
7.84437,
4.11822,
7.73243,
8.16779,
7.50725,
4.89209,
6.28632,
5.93133,
8.23422,
8.80662,
6.86181,
6.90161,
5.97109,
8.37274,
6.1324,
8.58223,
6.26041,
6.19714,
8.83858,
5.02823,
6.53406,
4.94321,
6.46434,
7.58531,
8.79829,
3.44372,
4.38396,
7.97783,
6.30135,
7.6139,
8.8632,
7.14381,
6.35142,
7.41854,
5.89967,
5.4361,
8.88114,
8.38241,
6.7143,
8.08667,
4.81073,
4.99441,
6.0604,
5.7585,
7.686,
5.72403,
6.68903,
8.51186,
7.21495,
5.58599,
8.77375,
6.99531,
4.62305,
5.45596,
8.71363,
5.21764,
6.72404,
8.50723,
7.66089,
7.2492,
6.1731,
6.28155,
5.25956,
8.76481,
5.28738,
6.80041,
5.00136,
6.27137,
4.88715,
5.66311,
8.96821,
7.62518,
4.49303,
6.8999,
6.18653,
7.62353,
5.26797,
6.30818,
8.75091,
5.22682,
6.91396,
8.83156,
8.97644,
4.98072,
5.22002,
8.44949,
3.64189,
7.70051,
5.454,
7.24937,
7.47875,
5.8002,
5.40274,
7.61586,
5.28606,
6.71455,
8.66638,
5.11625,
5.66604,
6.56109,
5.52685,
6.7965,
5.9041,
6.20023,
8.01596,
8.99811,
4.84864,
4.94429,
5.53183,
4.70004,
6.94536,
6.86479,
6.39941,
5.12868,
8.16441,
8.05361,
8.83382,
4.40875,
6.21299,
8.31721,
5.99746,
6.13926,
7.72945,
5.20223,
6.86095,
5.183,
7.51092,
8.49956,
7.68265,
8.99408,
6.40993,
6.04612,
4.12905,
7.04225,
4.33899,
5.71453,
8.10232,
6.69244,
8.63387,
5.67624,
4.64417,
6.84123,
5.9043,
4.71213,
8.23123,
5.00211,
8.42676,
6.81254,
4.11499,
6.12146,
5.77923,
6.70038,
4.52787,
5.7632,
5.59583,
6.60233,
5.57011,
7.64853,
3.37012,
5.84849,
6.5352,
5.7307,
4.2486,
8.55578,
4.60516,
6.04019,
8.47712,
4.00746,
6.04241,
8.44965,
8.19053,
6.63034,
7.3789,
4.62193,
7.26706,
8.46526,
8.48981,
5.91112,
5.68746,
7.58585,
4.60606,
5.96224,
4.33624,
5.201,
5.08792,
8.38858,
8.3854,
8.38379,
7.59093,
4.79026,
7.26037,
7.37631,
7.67865,
4.36201,
5.76338,
6.85426,
5.06256,
5.83644,
5.52457,
6.43461,
8.84871,
7.68169,
6.29525,
8.25434,
7.82436,
6.06282,
7.21737,
5.9913,
7.12784,
6.3329,
3.50612,
5.19803,
4.94444,
5.62464,
7.70534,
8.23105,
3.53071,
5.11078,
4.73921,
4.48016,
5.67041,
6.8633,
6.65612,
3.58703,
5.3655,
5.84459,
5.09844,
7.65193,
7.42143,
3.82056,
7.34648,
5.65678,
5.15114,
4.08664,
8.85835,
3.44579,
6.1396,
8.92349,
3.85085,
6.75439,
7.11673,
4.64145,
7.86186,
5.87164,
4.9815,
6.41565,
7.1668,
4.51993,
7.71981,
7.04416,
7.6527,
6.17844,
8.45957,
5.93233,
4.84919,
8.50099,
8.19291,
7.23766,
5.26005,
4.40513,
7.09172,
5.87765,
4.38964,
4.85278,
4.30482,
6.29605,
8.81498,
6.9329,
4.8081,
6.36249,
7.36317,
5.89809,
7.89598,
6.76941,
6.47239,
8.43861,
5.44945,
6.20295,
3.37149,
5.04378,
5.52549,
6.45649,
4.63402,
3.22653,
8.65684,
4.85636,
6.88472,
5.36066,
5.11308,
6.4047,
7.44259,
6.70223,
8.15972,
7.22989,
5.65507,
8.91146,
6.9378,
8.03705,
8.93738,
4.77778,
6.04027,
4.09842,
6.67132,
8.96107,
7.10758,
5.4704,
5.75726,
6.03449,
8.03455,
7.20312,
8.38266,
7.4456,
5.83184,
7.06892,
6.41179,
4.52211,
5.38736,
7.51541,
7.78534,
6.60505,
5.5876,
8.89239,
7.49174,
8.61059,
5.03924,
6.5323,
4.1597,
4.53097,
5.06776,
8.99583,
4.11686,
5.4276,
8.98056,
4.51286,
8.16593,
4.04629,
7.71885,
6.5108,
5.32329,
7.49895,
4.32715,
8.40041,
6.60146,
6.1728,
4.24057,
7.84756,
4.33488,
8.02943,
6.6436,
8.90289,
4.60036,
6.84769,
7.47611,
8.44158,
5.99604,
5.9653,
5.8115,
6.33175,
6.836,
6.76807,
8.13983,
5.34034,
8.81017,
5.49512,
5.15745,
6.95781,
8.94197,
8.65651,
6.38947,
8.41063,
7.32559,
5.0794,
5.64138,
8.49722,
7.28783,
5.08742,
6.78521,
8.11645,
4.0966,
6.9283,
5.95191,
6.91862,
5.67267,
4.66914,
7.79562,
7.88915,
3.47666,
6.48552,
5.69535,
8.03049,
8.80606,
6.25782,
7.57476,
4.02162,
6.23433,
7.66237,
7.92707,
6.22218,
7.08373,
6.35631,
6.21755,
5.02657,
7.81968,
8.79485,
5.79754,
7.65535,
7.09982,
7.15332,
5.73146,
5.4835,
4.69607,
8.40282,
8.86563,
6.14662,
7.49723,
7.83281,
5.64812,
6.74517,
5.5247,
4.86692,
6.90242,
5.56382,
4.91945,
8.78748,
8.91892,
8.0086,
7.36834,
5.55255,
6.15163,
4.70904,
5.5332,
8.87406,
5.91084,
8.97702,
8.9422,
4.54795,
7.59906,
6.16008,
6.2678,
4.79316,
5.766,
4.74259,
5.65983,
5.56641,
7.83453,
7.39732,
6.50318,
5.37484,
6.18223,
8.25643,
5.16514,
6.76341,
5.56466,
8.45027,
7.96694,
3.77071,
8.06529,
8.52489,
7.81787,
5.9646,
8.61096,
8.33811,
4.59511,
8.24258,
5.25415,
7.19029,
6.17983,
7.14333,
7.67227,
8.06726,
5.8942,
7.61427,
3.49898,
5.06289,
7.31791,
5.39542,
7.4956,
5.32236,
6.52822,
8.15125,
4.25369,
6.29676,
5.10226,
4.16865,
5.48507,
4.59742,
5.62444,
4.5249,
6.12301,
6.48564,
7.0461,
4.14299,
6.16497,
4.57273,
5.40557,
5.61805,
8.92726,
6.86283,
7.97776,
5.36381,
6.17184,
5.21335,
7.42788,
7.86201,
4.83528,
6.53465,
5.71023,
8.34906,
6.77614,
6.40499,
6.37239,
8.59818,
6.98013,
8.19941,
5.63077,
6.61975,
5.796,
6.98542,
5.8102,
8.63468,
4.11559,
5.94091,
6.72806,
4.97693,
5.4481,
8.89797,
4.10096,
8.10401,
5.47539,
8.61534,
4.36094,
5.54355,
5.58957,
6.76711,
8.11018,
8.6331,
6.23335,
6.12596,
8.19239,
5.04275,
6.83404,
7.03238,
7.28252,
5.32849,
4.86074,
6.54106,
6.05429,
7.22033,
8.69386,
3.77226,
5.54768,
5.32052,
5.63718,
5.76536,
4.6061,
4.67442,
7.72373,
6.5739,
6.55572,
8.15088,
4.31149,
5.92692,
8.427,
7.187,
4.8239,
5.42546,
7.42586,
7.35742,
4.57935,
8.18314,
7.53186,
5.22701,
7.75554,
4.4264,
6.91034,
8.90978,
7.0345,
4.42143,
6.14994,
5.90022,
6.86069,
8.66618,
7.14682,
8.10816,
5.20248,
4.58585,
7.53142,
6.00106,
6.28587,
5.88922,
7.96471,
8.49635,
7.84139,
5.23536,
4.46151,
8.91178,
5.80105,
6.11396,
3.85424,
7.83372,
6.74337,
6.38398,
6.11585,
5.11297,
8.60157,
3.86517,
4.91484,
5.37804,
3.76147,
6.07697,
6.56224,
8.94854,
5.87813,
4.75655,
4.91496,
5.15925,
7.59451,
7.26648,
5.36187,
6.08889,
5.0942,
5.52225,
5.9394,
6.5716,
5.30015,
7.06736,
6.9095,
4.61255,
4.68999,
7.21312,
4.17767;
}
