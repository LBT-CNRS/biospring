netcdf SpringNetwork {

dimensions:
	spatialdim = 3;
	particle_number = 183;
	particlename_length = 4;
	chainname_length = 4;
	resname_length = 4;

	springdim = 2; 
	spring_number = 1106;

variables:
	float   coordinates(particle_number, spatialdim); 
	        coordinates:units = "angstrom" ;
	        coordinates:long_name = "Particle coordinates";

	int     particleids(particle_number); 
	        particleids:long_name = "Particle ids in source database";

	char    particlenames(particle_number,particlename_length); 
	        particlenames:long_name = "Particle name";

	float   charges(particle_number);
	        charges:long_name = "Particle charge id";
	        charges:units = "electron" ;

	float   radii(particle_number);
	        radii:units = "A" ;
	        radii:long_name = "Particle radius";

	float   epsilon(particle_number);
	        epsilon:units = "kJ.mol-1" ;
	        epsilon:long_name = "Particle epsilon for Lennard-Jones";

	float   mass(particle_number);
	        mass:units = "Da" ;
	        mass:long_name = "Particle mass";

	float   surfaceaccessibility(particle_number);
	        surfaceaccessibility:units = "A2 or percent" ;
	        surfaceaccessibility:long_name = "Particle surface accessibility";

	float   hydrophobicityscale(particle_number);
	        hydrophobicityscale:units = "kJ.mol-1" ;
	        hydrophobicityscale:long_name = "Particle hydrophobicity scale (transfer energy)";

	char    resnames(particle_number,resname_length); 
	        resnames:long_name = "particle residue name";

	int     resids(particle_number); 
	        resids:long_name = "particle residue id";

	char    chainnames(particle_number,chainname_length); 
	        chainnames:long_name = "Chain name ";

	byte    dynamicstate(particle_number); 
	        dynamicstate:long_name = "particle dynamic state (static 0 or dynamic 1)";

	int     springs(spring_number,springdim); 
	        springs:long_name = "Spring between particle referenced by 2 particle ids"; 

	float   springsstiffness(spring_number); 
	        springsstiffness:long_name = "Spring stiffness";
	float   springsequilibrium(spring_number); 
	        springsequilibrium:long_name = "Spring distance equilibrium";
data:
	particleids = 
1,
2,
3,
4,
5,
6,
7,
8,
9,
10,
11,
12,
13,
14,
15,
16,
17,
18,
19,
20,
21,
22,
23,
24,
25,
26,
27,
28,
29,
30,
31,
32,
33,
34,
35,
36,
37,
38,
39,
40,
41,
42,
43,
44,
45,
46,
47,
48,
49,
50,
51,
52,
53,
54,
55,
56,
57,
58,
59,
60,
61,
62,
63,
64,
65,
66,
67,
68,
69,
70,
71,
72,
73,
74,
75,
76,
77,
78,
79,
80,
81,
82,
83,
84,
85,
86,
87,
88,
89,
90,
91,
92,
93,
94,
95,
96,
97,
98,
99,
100,
101,
102,
103,
104,
105,
106,
107,
108,
109,
110,
111,
112,
113,
114,
115,
116,
117,
118,
119,
120,
121,
122,
123,
124,
125,
126,
127,
128,
129,
130,
131,
132,
133,
134,
135,
136,
137,
138,
139,
140,
141,
142,
143,
144,
145,
146,
147,
148,
149,
150,
151,
152,
153,
154,
155,
156,
157,
158,
159,
160,
161,
162,
163,
164,
165,
166,
167,
168,
169,
170,
171,
172,
173,
174,
175,
176,
177,
178,
179,
180,
181,
182,
183;
	coordinates = 
9.27257, 34.0063, 15.0073,
10.826, 29.9498, 14.937,
14.3379, 32.3195, 12.3651,
16.3871, 27.5676, 14.4209,
19.985, 30.2409, 15.4413,
22.8017, 26.984, 14.4686,
25.7259, 30.35, 16.929,
29.0214, 28.97, 15.128,
32.6787, 29.158, 14.972,
35.7699, 30.3063, 15.2976,
37.514, 29.1342, 18.69,
37.6656, 32.2484, 20.7806,
34.8493, 34.0841, 18.1909,
32.578, 34.8545, 21.299,
30.101, 30.8927, 20.5457,
29.3092, 32.7348, 24.6374,
29.6876, 36.4533, 24.94,
26.8071, 36.4533, 21.56,
24.7861, 32.9681, 23.414,
25.5082, 35.9865, 28.7448,
23.2475, 38.6895, 24.775,
20.9878, 36.4891, 22.1399,
19.7917, 32.6722, 27.1954,
20.6584, 38.6414, 28.7202,
19.4335, 41.9021, 24.6698,
15.2835, 37.0991, 23.416,
13.2723, 36.6217, 27.4599,
10.8032, 33.7516, 24.4406,
15.2975, 32.2915, 23.3545,
14.6393, 26.7528, 23.1978,
19.9474, 27.5401, 24.843,
19.3334, 24.1284, 23.3296,
19.8884, 22.7739, 27.0603,
22.0994, 19.64, 26.2676,
21.987, 16.196, 26.5436,
24.3407, 14.5151, 29.4147,
25.497, 10.518, 29.6977,
27.4255, 14.8075, 33.3431,
26.226, 12.9474, 36.4524,
24.725, 15.4484, 38.2364,
29.1182, 19.298, 37.3449,
27.4427, 19.4937, 42.8023,
23.5243, 21.784, 41.8913,
24.2172, 20.6993, 37.8339,
19.1669, 21.8646, 37.5831,
17.2479, 18.3076, 34.7534,
17.4062, 21.3492, 31.9397,
18.6823, 24.3683, 33.583,
22.5823, 23.057, 33.7578,
24.0567, 19.7922, 30.4262,
18.1955, 17.8503, 29.2456,
21.4328, 15.6383, 33.749,
19.7389, 11.1942, 29.8776,
20.6864, 6.34675, 30.8195,
23.5844, 5.986, 28.9946,
20.8526, 3.17443, 27.0321,
16.2348, 7.46782, 26.2682,
22.1576, 9.95064, 24.3092,
22.291, 4.88578, 21.5724,
17.3317, 4.114, 22.9983,
17.1339, 9.19937, 21.6706,
21.2996, 8.24675, 18.5569,
19.1558, 4.5695, 17.1185,
14.5572, 6.86144, 18.0778,
16.4615, 10.7615, 15.6343,
14.6976, 12.0587, 18.5444,
19.934, 13.3175, 18.9741,
19.4709, 17.3528, 15.8631,
24.2418, 17.1602, 17.7352,
26.5438, 11.739, 18.8669,
29.2836, 13.9096, 21.0648,
31.7813, 10.6176, 22.3879,
32.4225, 14.2346, 25.783,
35.909, 14.4347, 28.665,
36.9148, 10.1092, 25.2603,
33.9762, 8.676, 26.078,
33.9318, 9.47462, 30.2506,
30.5587, 12.3059, 28.9038,
27.7259, 9.50909, 24.361,
26.5276, 15.0642, 24.4042,
23.447, 16.6658, 22.833,
21.0453, 18.6999, 20.3523,
17.4164, 16.777, 22.4726,
14.7554, 17.3402, 18.7554,
11.6397, 16.0254, 21.4696,
13.083, 20.4594, 22.5664,
13.899, 22.3554, 18.7237,
10.9535, 20.2382, 15.1923,
8.2396, 22.4366, 20.148,
9.5892, 25.6502, 19.7682,
9.0538, 25.8148, 16.2822,
5.6428, 24.7654, 16.6436,
5.06357, 27.0519, 19.6491,
6.85775, 30.1823, 17.7302,
9.18143, 30.0831, 20.2727,
12.5033, 31.8569, 19.4676,
15.549, 28.4306, 18.7414,
20.0191, 29.782, 20.4755,
21.3995, 25.7996, 18.843,
26.3921, 27.0797, 21.7803,
27.2724, 24.0217, 18.1213,
30.9526, 22.227, 16.4964,
31.7725, 23.9569, 12.6406,
30.0242, 19.51, 13.176,
27.0127, 20.1832, 14.5343,
26.0454, 22.549, 12.565,
28.0243, 20.2261, 8.15764,
24.2486, 17.8532, 11.6352,
21.655, 20.5879, 13.2451,
21.1074, 22.2953, 7.77422,
22.4226, 16.6264, 7.394,
18.3236, 16.7671, 11.1887,
15.9396, 21.2014, 11.4085,
16.7347, 21.4827, 6.95671,
13.8909, 23.772, 8.85944,
17.7322, 25.7674, 10.1356,
19.7729, 29.259, 10.2657,
23.8683, 27.9254, 9.84943,
25.1039, 31.6296, 12.2817,
30.915, 31.6185, 10.9344,
30.573, 34.5412, 15.1699,
33.402, 36.3244, 12.8036,
36.6611, 37.3569, 13.4354,
37.4493, 41.2742, 13.8906,
40.502, 39.976, 12.389,
44.1064, 35.1571, 11.8332,
46.2171, 40.6596, 13.5792,
42.0645, 40.0154, 17.1658,
41.5218, 35.2044, 16.6691,
46.9572, 35.4206, 15.5557,
46.434, 37.5302, 19.5506,
41.9072, 36.9629, 21.0205,
44.5199, 32.1248, 20.1539,
49.1802, 34.06, 21.2559,
48.266, 35.6332, 24.5585,
49.5555, 37.9561, 28.3077,
52.6345, 33.1087, 26.0245,
51.95, 31.2531, 28.9109,
50.2699, 27.7196, 25.6978,
53.8353, 25.7527, 24.4676,
54.4046, 27.35, 20.6594,
53.2773, 23.0706, 19.7156,
49.8296, 24.245, 21.6901,
49.9959, 28.6246, 20.3859,
51.0624, 27.0277, 15.5391,
46.5178, 21.7872, 18.1956,
44.9608, 26.7786, 20.4908,
46.9474, 29.5276, 15.096,
45.9125, 24.8289, 12.1709,
42.3983, 24.7829, 14.3124,
41.5082, 28.6544, 13.2942,
44.2276, 30.3499, 8.71455,
40.6845, 24.6595, 9.6415,
37.553, 26.8542, 12.9288,
38.0903, 30.9819, 9.60213,
36.9848, 27.9116, 5.9996,
33.395, 27.2694, 6.9644,
33.0622, 31.8202, 6.33556,
30.5993, 29.5665, 3.06375,
28.7676, 25.803, 4.09825,
27.8394, 28.261, 8.14382,
23.0222, 29.6459, 6.067,
23.2497, 34.0417, 7.33022,
28.1223, 35.6089, 8.39,
27.9454, 37.7721, 12.2477,
31.4313, 40.4811, 12.0044,
32.3047, 39.8986, 17.0999,
33.4888, 44.3316, 13.4081,
31.1475, 46.3913, 20.737,
29.1469, 41.7795, 22.1991,
27.2734, 45.129, 22.5544,
26.2132, 44.7436, 17.7092,
26.4636, 41.2746, 17.0808,
23.6752, 40.6985, 19.6947,
21.6726, 43.0094, 17.5042,
23.4756, 41.5076, 13.1856,
21.9166, 37.374, 15.8504,
17.976, 40.0223, 17.6967,
17.1954, 40.4922, 13.6594,
18.0501, 36.2669, 12.3044,
16.2684, 35.1711, 16.4154,
12.8297, 38.3559, 16.5859,
13.6722, 41.3877, 13.838;
	charges = 
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
1,
0,
0,
1,
-1,
1,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
1,
0,
0,
-1,
0,
-1,
0,
0,
-1,
0,
1,
0,
0,
-1,
0,
0,
1,
0,
0,
0,
0,
0,
-1,
0,
0,
-1,
0,
0,
-1,
0,
0,
-1,
0,
1,
0,
0,
0,
1,
1,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
-1,
0,
0,
0,
0,
1,
0,
0,
1,
1,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
1,
0,
0,
0,
1,
0,
0,
-1,
0,
0,
-1,
0,
0,
0,
1,
1,
0,
-1,
0,
0,
1,
0,
-1,
0,
0,
0,
0,
0,
-1,
0,
-1,
1,
0,
0,
0,
0,
1,
1,
0,
-1,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0;
	radii = 
3.3,
2.58,
3.47,
3.3,
3.3,
3.3,
3.49,
2.89,
2.58,
3.2,
2.89,
2.88,
3.3,
2.58,
3.44,
2.89,
3.12,
3.3,
3.3,
3.47,
3.03,
3.49,
3.47,
3.22,
3.47,
3.47,
3.2,
3.13,
3.49,
3.38,
3.64,
2.89,
3.3,
2.89,
2.88,
3.12,
3.12,
3.47,
2.88,
3.2,
3.47,
3.2,
2.58,
3.22,
3.3,
3,
2.58,
3.3,
3,
3.66,
3.38,
3.64,
3.47,
3,
3.2,
3.12,
3.47,
3.64,
3.34,
3.34,
3.49,
3.47,
3,
3.34,
2.58,
3.22,
3.49,
3.49,
3.22,
3.85,
2.88,
3.22,
3.47,
3.38,
2.58,
2.58,
3.49,
3.38,
3.47,
2.89,
2.58,
3.12,
3.49,
2.88,
3.34,
3.2,
3.3,
3.47,
2.88,
2.88,
2.88,
2.88,
3.12,
2.58,
3.3,
3.2,
3.3,
3.49,
3.47,
3.22,
3.3,
3,
3.49,
2.88,
2.58,
2.88,
3.47,
2.88,
3.47,
3.44,
3.44,
3.12,
3.47,
3.2,
3.22,
2.88,
3.3,
3.12,
3.3,
3.64,
3.49,
2.88,
3.2,
3.2,
2.89,
3.85,
3.34,
3,
3.49,
3.34,
2.88,
3.47,
3.49,
3.47,
2.58,
3.47,
2.58,
3.12,
3.22,
3.12,
2.88,
3,
3.3,
3.47,
3.34,
3.47,
3.47,
3.49,
3,
3.12,
2.88,
3.47,
3.47,
3.22,
3.49,
2.88,
2.88,
3.34,
2.58,
3,
3.64,
3,
3.44,
3.3,
3.3,
3.3,
3.13,
3.47,
3.47,
3.49,
3.22,
2.89,
2.88,
3.03,
2.88,
3.22,
3.49,
3.3,
2.89,
3.49,
3.49,
3.3,
2.58;
	epsilon = 
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1;
	mass = 
117,
75,
174,
117,
117,
117,
131,
105,
75,
115,
105,
89,
117,
75,
146,
105,
119,
117,
117,
174,
121,
131,
174,
147,
174,
131,
115,
132,
131,
155,
165,
105,
117,
105,
89,
119,
119,
174,
89,
115,
174,
115,
75,
147,
117,
133,
75,
117,
133,
181,
155,
165,
131,
133,
115,
119,
174,
165,
146,
146,
131,
131,
133,
146,
75,
147,
131,
131,
147,
204,
89,
147,
131,
155,
75,
75,
131,
155,
174,
105,
75,
119,
131,
89,
146,
115,
117,
174,
89,
89,
89,
89,
119,
75,
117,
115,
117,
131,
131,
147,
117,
133,
131,
89,
75,
89,
174,
89,
131,
146,
146,
119,
149,
115,
147,
89,
117,
119,
117,
165,
131,
89,
115,
115,
105,
204,
146,
133,
131,
146,
89,
174,
131,
131,
75,
174,
75,
119,
147,
119,
89,
133,
117,
131,
146,
174,
174,
131,
133,
119,
89,
174,
131,
147,
131,
89,
89,
146,
75,
133,
165,
133,
146,
117,
117,
117,
132,
174,
174,
131,
147,
105,
89,
121,
89,
147,
131,
117,
105,
131,
131,
117,
75;
	surfaceaccessibility = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	hydrophobicityscale = 
5.04836,
0,
-4.17938,
5.04836,
5.04836,
5.04836,
7.0346,
-0.16552,
0,
2.97936,
-0.16552,
1.28278,
5.04836,
0,
-4.09662,
-0.16552,
1.07588,
5.04836,
5.04836,
-4.17938,
6.37252,
7.0346,
-4.17938,
-2.64832,
-4.17938,
7.4484,
2.97936,
-2.4828,
7.0346,
0.53794,
7.40702,
-0.16552,
5.04836,
-0.16552,
1.28278,
1.07588,
1.07588,
-4.17938,
1.28278,
2.97936,
-4.17938,
2.97936,
0,
-2.64832,
5.04836,
-3.18626,
0,
5.04836,
-3.18626,
3.97248,
0.53794,
7.40702,
7.4484,
-3.18626,
2.97936,
1.07588,
-4.17938,
7.40702,
-0.91036,
-0.91036,
7.0346,
7.4484,
-3.18626,
-0.91036,
0,
-2.64832,
7.0346,
7.0346,
-2.64832,
9.3105,
1.28278,
-2.64832,
7.4484,
0.53794,
0,
0,
7.0346,
0.53794,
-4.17938,
-0.16552,
0,
1.07588,
7.0346,
1.28278,
-0.91036,
2.97936,
5.04836,
-4.17938,
1.28278,
1.28278,
1.28278,
1.28278,
1.07588,
0,
5.04836,
2.97936,
5.04836,
7.0346,
7.4484,
-2.64832,
5.04836,
-3.18626,
7.0346,
1.28278,
0,
1.28278,
-4.17938,
1.28278,
7.4484,
-4.09662,
-4.09662,
1.07588,
5.08974,
2.97936,
-2.64832,
1.28278,
5.04836,
1.07588,
5.04836,
7.40702,
7.0346,
1.28278,
2.97936,
2.97936,
-0.16552,
9.3105,
-0.91036,
-3.18626,
7.0346,
-0.91036,
1.28278,
-4.17938,
7.0346,
7.4484,
0,
-4.17938,
0,
1.07588,
-2.64832,
1.07588,
1.28278,
-3.18626,
5.04836,
7.4484,
-0.91036,
-4.17938,
-4.17938,
7.0346,
-3.18626,
1.07588,
1.28278,
-4.17938,
7.4484,
-2.64832,
7.0346,
1.28278,
1.28278,
-0.91036,
0,
-3.18626,
7.40702,
-3.18626,
-4.09662,
5.04836,
5.04836,
5.04836,
-2.4828,
-4.17938,
-4.17938,
7.0346,
-2.64832,
-0.16552,
1.28278,
6.37252,
1.28278,
-2.64832,
7.0346,
5.04836,
-0.16552,
7.0346,
7.0346,
5.04836,
0;
	particlenames = 
"VCA",
"GCA",
"RCA",
"VCA",
"VCA",
"VCA",
"LCA",
"SCA",
"GCA",
"PCA",
"SCA",
"ACA",
"VCA",
"GCA",
"KCA",
"SCA",
"TCA",
"VCA",
"VCA",
"RCA",
"CCA",
"LCA",
"RCA",
"ECA",
"RCA",
"ICA",
"PCA",
"NCA",
"LCA",
"HCA",
"FCA",
"SCA",
"VCA",
"SCA",
"ACA",
"TCA",
"TCA",
"RCA",
"ACA",
"PCA",
"RCA",
"PCA",
"GCA",
"ECA",
"VCA",
"DCA",
"GCA",
"VCA",
"DCA",
"YCA",
"HCA",
"FCA",
"ICA",
"DCA",
"PCA",
"TCA",
"RCA",
"FCA",
"QCA",
"QCA",
"LCA",
"ICA",
"DCA",
"QCA",
"GCA",
"ECA",
"LCA",
"LCA",
"ECA",
"WCA",
"ACA",
"ECA",
"ICA",
"HCA",
"GCA",
"GCA",
"LCA",
"HCA",
"RCA",
"SCA",
"GCA",
"TCA",
"LCA",
"ACA",
"QCA",
"PCA",
"VCA",
"RCA",
"ACA",
"ACA",
"ACA",
"ACA",
"TCA",
"GCA",
"VCA",
"PCA",
"VCA",
"LCA",
"ICA",
"ECA",
"VCA",
"DCA",
"LCA",
"ACA",
"GCA",
"ACA",
"RCA",
"ACA",
"ICA",
"KCA",
"KCA",
"TCA",
"MCA",
"PCA",
"ECA",
"ACA",
"VCA",
"TCA",
"VCA",
"FCA",
"LCA",
"ACA",
"PCA",
"PCA",
"SCA",
"WCA",
"QCA",
"DCA",
"LCA",
"QCA",
"ACA",
"RCA",
"LCA",
"ICA",
"GCA",
"RCA",
"GCA",
"TCA",
"ECA",
"TCA",
"ACA",
"DCA",
"VCA",
"ICA",
"QCA",
"RCA",
"RCA",
"LCA",
"DCA",
"TCA",
"ACA",
"RCA",
"ICA",
"ECA",
"LCA",
"ACA",
"ACA",
"QCA",
"GCA",
"DCA",
"FCA",
"DCA",
"KCA",
"VCA",
"VCA",
"VCA",
"NCA",
"RCA",
"RCA",
"LCA",
"ECA",
"SCA",
"ACA",
"CCA",
"ACA",
"ECA",
"LCA",
"VCA",
"SCA",
"LCA",
"LCA",
"VCA",
"GCA";
	resnames = 
"VAL",
"GLY",
"ARG",
"VAL",
"VAL",
"VAL",
"LEU",
"SER",
"GLY",
"PRO",
"SER",
"ALA",
"VAL",
"GLY",
"LYS",
"SER",
"THR",
"VAL",
"VAL",
"ARG",
"CYS",
"LEU",
"ARG",
"GLU",
"ARG",
"ILE",
"PRO",
"ASN",
"LEU",
"HIS",
"PHE",
"SER",
"VAL",
"SER",
"ALA",
"THR",
"THR",
"ARG",
"ALA",
"PRO",
"ARG",
"PRO",
"GLY",
"GLU",
"VAL",
"ASP",
"GLY",
"VAL",
"ASP",
"TYR",
"HIS",
"PHE",
"ILE",
"ASP",
"PRO",
"THR",
"ARG",
"PHE",
"GLN",
"GLN",
"LEU",
"ILE",
"ASP",
"GLN",
"GLY",
"GLU",
"LEU",
"LEU",
"GLU",
"TRP",
"ALA",
"GLU",
"ILE",
"HIS",
"GLY",
"GLY",
"LEU",
"HIS",
"ARG",
"SER",
"GLY",
"THR",
"LEU",
"ALA",
"GLN",
"PRO",
"VAL",
"ARG",
"ALA",
"ALA",
"ALA",
"ALA",
"THR",
"GLY",
"VAL",
"PRO",
"VAL",
"LEU",
"ILE",
"GLU",
"VAL",
"ASP",
"LEU",
"ALA",
"GLY",
"ALA",
"ARG",
"ALA",
"ILE",
"LYS",
"LYS",
"THR",
"MET",
"PRO",
"GLU",
"ALA",
"VAL",
"THR",
"VAL",
"PHE",
"LEU",
"ALA",
"PRO",
"PRO",
"SER",
"TRP",
"GLN",
"ASP",
"LEU",
"GLN",
"ALA",
"ARG",
"LEU",
"ILE",
"GLY",
"ARG",
"GLY",
"THR",
"GLU",
"THR",
"ALA",
"ASP",
"VAL",
"ILE",
"GLN",
"ARG",
"ARG",
"LEU",
"ASP",
"THR",
"ALA",
"ARG",
"ILE",
"GLU",
"LEU",
"ALA",
"ALA",
"GLN",
"GLY",
"ASP",
"PHE",
"ASP",
"LYS",
"VAL",
"VAL",
"VAL",
"ASN",
"ARG",
"ARG",
"LEU",
"GLU",
"SER",
"ALA",
"CYS",
"ALA",
"GLU",
"LEU",
"VAL",
"SER",
"LEU",
"LEU",
"VAL",
"GLY";
	resids = 
1,
2,
3,
4,
5,
6,
7,
8,
9,
10,
11,
12,
13,
14,
15,
16,
17,
18,
19,
20,
21,
22,
23,
24,
25,
26,
27,
28,
29,
30,
31,
32,
33,
34,
35,
36,
37,
38,
39,
40,
41,
42,
43,
44,
45,
46,
47,
48,
49,
50,
51,
52,
53,
54,
55,
56,
57,
58,
59,
60,
61,
62,
63,
64,
65,
66,
67,
68,
69,
70,
71,
72,
73,
74,
75,
76,
77,
78,
79,
80,
81,
82,
83,
84,
85,
86,
87,
88,
89,
90,
91,
92,
93,
94,
95,
96,
97,
98,
99,
100,
101,
102,
103,
104,
105,
106,
107,
108,
109,
110,
111,
112,
113,
114,
115,
116,
117,
118,
119,
120,
121,
122,
123,
124,
125,
126,
127,
128,
129,
130,
131,
132,
133,
134,
135,
136,
137,
138,
139,
140,
141,
142,
143,
144,
145,
146,
147,
148,
149,
150,
151,
152,
153,
154,
155,
156,
157,
158,
159,
160,
161,
162,
163,
164,
165,
166,
167,
168,
169,
170,
171,
172,
173,
174,
175,
176,
177,
178,
179,
180,
181,
182,
183;
	chainnames = 
"1",
"2",
"3",
"4",
"5",
"6",
"7",
"8",
"9",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"2",
"2",
"2",
"2",
"2",
"2",
"2",
"2",
"2",
"2",
"3",
"3",
"3",
"3",
"3",
"3",
"3",
"3",
"3",
"3",
"4",
"4",
"4",
"4",
"4",
"4",
"4",
"4",
"4",
"4",
"5",
"5",
"5",
"5",
"5",
"5",
"5",
"5",
"5",
"5",
"6",
"6",
"6",
"6",
"6",
"6",
"6",
"6",
"6",
"6",
"7",
"7",
"7",
"7",
"7",
"7",
"7",
"7",
"7",
"7",
"8",
"8",
"8",
"8",
"8",
"8",
"8",
"8",
"8",
"8",
"9",
"9",
"9",
"9",
"9",
"9",
"9",
"9",
"9",
"9",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1",
"1";
	dynamicstate = 
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1;
	springs = 
0, 1,
0, 2,
0, 180,
0, 181,
0, 182,
0, 90,
0, 93,
0, 94,
0, 95,
1, 2,
1, 3,
1, 180,
1, 181,
1, 89,
1, 90,
1, 91,
1, 92,
1, 93,
1, 94,
1, 95,
1, 96,
2, 3,
2, 4,
2, 115,
2, 116,
2, 178,
2, 179,
2, 180,
2, 181,
2, 95,
2, 96,
3, 97,
3, 98,
3, 4,
3, 5,
3, 108,
3, 112,
3, 114,
3, 115,
3, 116,
3, 117,
3, 29,
3, 180,
3, 86,
3, 89,
3, 90,
3, 95,
3, 96,
4, 97,
4, 98,
4, 5,
4, 6,
4, 115,
4, 116,
4, 117,
4, 118,
4, 176,
4, 179,
4, 180,
4, 95,
4, 96,
5, 97,
5, 98,
5, 99,
5, 100,
5, 6,
5, 104,
5, 7,
5, 105,
5, 108,
5, 109,
5, 115,
5, 116,
5, 117,
5, 118,
5, 160,
5, 161,
5, 96,
6, 97,
6, 98,
6, 99,
6, 100,
6, 7,
6, 105,
6, 8,
6, 14,
6, 15,
6, 17,
6, 18,
6, 117,
6, 118,
6, 119,
6, 120,
6, 176,
7, 99,
7, 100,
7, 101,
7, 102,
7, 105,
7, 8,
7, 9,
7, 12,
7, 14,
7, 117,
7, 118,
7, 119,
7, 120,
7, 121,
7, 160,
8, 100,
8, 101,
8, 102,
8, 9,
8, 10,
8, 11,
8, 12,
8, 13,
8, 14,
8, 118,
8, 119,
8, 120,
8, 121,
8, 153,
8, 154,
8, 156,
8, 160,
9, 102,
9, 10,
9, 11,
9, 12,
9, 13,
9, 14,
9, 119,
9, 120,
9, 121,
9, 122,
9, 128,
9, 149,
9, 150,
9, 153,
9, 154,
10, 11,
10, 12,
10, 13,
10, 14,
10, 128,
10, 132,
10, 146,
10, 149,
10, 150,
10, 153,
11, 12,
11, 13,
11, 14,
11, 128,
11, 131,
11, 132,
12, 13,
12, 14,
12, 15,
12, 16,
12, 119,
12, 120,
12, 121,
12, 122,
12, 123,
12, 128,
12, 131,
12, 166,
13, 14,
13, 15,
13, 16,
13, 17,
13, 18,
13, 120,
13, 121,
13, 166,
13, 169,
14, 99,
14, 100,
14, 15,
14, 16,
14, 17,
14, 18,
14, 120,
15, 99,
15, 16,
15, 17,
15, 18,
15, 19,
15, 20,
16, 17,
16, 18,
16, 19,
16, 20,
16, 166,
16, 169,
17, 18,
17, 19,
17, 20,
17, 21,
17, 120,
17, 166,
17, 169,
17, 170,
17, 172,
17, 173,
17, 176,
18, 97,
18, 99,
18, 19,
18, 20,
18, 21,
18, 22,
18, 23,
18, 30,
18, 173,
19, 20,
19, 21,
19, 22,
19, 23,
20, 21,
20, 22,
20, 23,
20, 24,
20, 25,
20, 169,
20, 170,
20, 172,
20, 173,
20, 174,
20, 177,
21, 97,
21, 22,
21, 23,
21, 24,
21, 25,
21, 28,
21, 172,
21, 173,
21, 174,
21, 176,
21, 177,
21, 180,
22, 97,
22, 23,
22, 25,
22, 26,
22, 28,
22, 29,
22, 30,
23, 24,
23, 25,
23, 26,
24, 25,
24, 26,
24, 170,
24, 173,
24, 174,
24, 177,
25, 95,
25, 26,
25, 27,
25, 28,
25, 177,
25, 180,
25, 181,
26, 27,
26, 28,
27, 28,
27, 29,
27, 93,
27, 94,
27, 95,
28, 97,
28, 29,
28, 30,
28, 180,
28, 94,
28, 95,
28, 96,
29, 97,
29, 98,
29, 30,
29, 31,
29, 32,
29, 85,
29, 86,
29, 88,
29, 89,
29, 90,
29, 94,
29, 95,
29, 96,
30, 97,
30, 98,
30, 99,
30, 31,
30, 32,
30, 33,
30, 96,
31, 97,
31, 98,
31, 99,
31, 32,
31, 33,
31, 34,
31, 50,
31, 80,
31, 81,
31, 82,
31, 85,
31, 86,
31, 96,
32, 98,
32, 33,
32, 34,
32, 46,
32, 47,
32, 48,
32, 49,
32, 50,
32, 80,
32, 81,
32, 82,
32, 85,
33, 34,
33, 35,
33, 46,
33, 48,
33, 49,
33, 50,
33, 51,
33, 79,
33, 80,
33, 81,
33, 82,
34, 35,
34, 36,
34, 37,
34, 46,
34, 49,
34, 50,
34, 51,
34, 52,
34, 57,
34, 66,
34, 79,
34, 80,
34, 81,
34, 82,
35, 49,
35, 50,
35, 51,
35, 52,
35, 54,
35, 57,
35, 72,
35, 77,
35, 78,
35, 79,
35, 80,
35, 36,
35, 37,
35, 38,
35, 39,
36, 51,
36, 52,
36, 53,
36, 54,
36, 57,
36, 72,
36, 76,
36, 77,
36, 78,
36, 79,
36, 37,
36, 38,
37, 49,
37, 51,
37, 76,
37, 77,
37, 79,
37, 38,
37, 39,
37, 40,
37, 43,
38, 51,
38, 77,
38, 39,
38, 40,
38, 43,
39, 49,
39, 51,
39, 40,
39, 41,
39, 42,
39, 43,
39, 44,
39, 45,
40, 48,
40, 49,
40, 41,
40, 42,
40, 43,
41, 42,
41, 43,
42, 48,
42, 43,
42, 44,
43, 47,
43, 48,
43, 49,
43, 51,
43, 44,
43, 45,
44, 45,
44, 46,
44, 47,
44, 48,
44, 49,
44, 51,
45, 47,
45, 48,
45, 49,
45, 50,
45, 51,
45, 52,
45, 46,
46, 47,
46, 48,
46, 49,
46, 50,
46, 51,
47, 48,
47, 49,
47, 50,
48, 49,
48, 50,
48, 51,
49, 50,
49, 51,
49, 79,
49, 80,
50, 51,
50, 52,
50, 80,
50, 82,
50, 85,
51, 52,
52, 53,
52, 54,
52, 55,
52, 56,
52, 57,
52, 60,
53, 54,
53, 55,
53, 56,
53, 57,
53, 59,
54, 55,
54, 56,
54, 57,
54, 58,
54, 59,
54, 78,
55, 56,
55, 57,
55, 58,
55, 59,
55, 60,
56, 57,
56, 58,
56, 59,
56, 60,
56, 63,
57, 58,
57, 59,
57, 60,
57, 61,
57, 66,
57, 69,
57, 70,
57, 78,
57, 79,
57, 80,
57, 82,
58, 59,
58, 60,
58, 61,
58, 62,
58, 63,
58, 69,
58, 78,
59, 60,
59, 61,
59, 62,
59, 63,
60, 61,
60, 62,
60, 63,
60, 64,
60, 65,
60, 66,
60, 82,
60, 83,
60, 84,
61, 62,
61, 63,
61, 64,
61, 65,
61, 66,
61, 69,
61, 78,
62, 63,
62, 64,
62, 65,
62, 66,
63, 64,
63, 65,
63, 66,
64, 111,
64, 65,
64, 66,
64, 67,
64, 83,
65, 66,
65, 67,
65, 82,
65, 83,
65, 84,
66, 111,
66, 67,
66, 68,
66, 69,
66, 79,
66, 80,
66, 81,
66, 82,
66, 83,
67, 104,
67, 107,
67, 108,
67, 110,
67, 111,
67, 112,
67, 68,
67, 80,
67, 81,
67, 82,
67, 83,
67, 86,
68, 100,
68, 101,
68, 103,
68, 104,
68, 105,
68, 107,
68, 108,
68, 111,
68, 69,
68, 70,
68, 79,
68, 80,
68, 81,
68, 82,
69, 70,
69, 71,
69, 78,
69, 79,
69, 80,
69, 81,
70, 71,
70, 72,
70, 75,
70, 77,
70, 78,
70, 79,
70, 80,
71, 72,
71, 73,
71, 74,
71, 75,
71, 76,
71, 77,
71, 78,
71, 79,
72, 73,
72, 74,
72, 75,
72, 76,
72, 77,
72, 78,
72, 79,
73, 74,
73, 75,
73, 76,
73, 77,
74, 75,
74, 76,
74, 77,
75, 76,
75, 77,
75, 78,
76, 77,
76, 78,
77, 78,
77, 79,
78, 79,
78, 80,
79, 80,
79, 81,
80, 81,
80, 82,
81, 98,
81, 100,
81, 104,
81, 108,
81, 82,
81, 83,
81, 85,
81, 86,
82, 83,
82, 84,
82, 85,
82, 86,
83, 111,
83, 112,
83, 84,
83, 85,
83, 86,
83, 87,
83, 88,
84, 85,
84, 86,
84, 87,
84, 88,
85, 86,
85, 87,
85, 88,
85, 89,
86, 98,
86, 112,
86, 87,
86, 88,
86, 89,
86, 90,
86, 91,
86, 96,
87, 112,
87, 114,
87, 88,
87, 89,
87, 90,
87, 91,
88, 94,
88, 89,
88, 90,
88, 91,
88, 92,
88, 93,
89, 90,
89, 91,
89, 92,
89, 93,
89, 94,
89, 95,
89, 96,
90, 91,
90, 92,
90, 93,
90, 94,
90, 95,
90, 96,
91, 94,
91, 92,
91, 93,
92, 94,
92, 95,
92, 93,
93, 94,
93, 95,
93, 96,
94, 95,
94, 96,
95, 97,
95, 180,
95, 181,
95, 96,
96, 97,
96, 98,
96, 180,
97, 98,
97, 99,
97, 180,
98, 99,
98, 100,
98, 105,
98, 108,
99, 100,
99, 101,
100, 101,
100, 102,
100, 103,
100, 104,
100, 105,
100, 108,
101, 102,
101, 103,
101, 104,
101, 105,
101, 153,
102, 103,
102, 104,
102, 105,
102, 106,
102, 119,
102, 153,
102, 156,
102, 160,
103, 104,
103, 105,
103, 106,
103, 107,
103, 108,
104, 105,
104, 106,
104, 107,
104, 108,
105, 106,
105, 107,
105, 108,
105, 109,
105, 110,
105, 117,
105, 160,
106, 107,
106, 108,
106, 156,
106, 109,
106, 110,
106, 159,
106, 160,
106, 117,
107, 108,
107, 109,
107, 110,
107, 111,
107, 112,
108, 109,
108, 110,
108, 111,
108, 112,
108, 113,
108, 115,
108, 117,
109, 110,
109, 111,
109, 112,
109, 113,
109, 114,
109, 115,
109, 116,
109, 117,
109, 161,
110, 111,
110, 112,
110, 113,
111, 112,
111, 113,
111, 114,
112, 113,
112, 114,
112, 115,
112, 116,
113, 114,
113, 115,
113, 116,
114, 115,
114, 116,
115, 161,
115, 116,
115, 117,
116, 117,
116, 118,
116, 160,
116, 161,
116, 162,
116, 179,
117, 118,
117, 119,
117, 159,
117, 160,
117, 161,
117, 162,
117, 163,
118, 119,
118, 120,
118, 160,
118, 161,
118, 162,
118, 163,
118, 164,
118, 176,
118, 179,
119, 120,
119, 121,
119, 122,
119, 153,
119, 154,
119, 155,
119, 156,
119, 157,
119, 158,
119, 160,
119, 162,
119, 163,
119, 164,
119, 165,
120, 121,
120, 122,
120, 163,
120, 164,
120, 165,
120, 166,
120, 172,
121, 122,
121, 123,
121, 124,
121, 154,
121, 157,
121, 163,
121, 164,
121, 165,
121, 166,
121, 167,
122, 123,
122, 124,
122, 125,
122, 127,
122, 128,
122, 154,
122, 164,
122, 165,
122, 166,
122, 167,
123, 124,
123, 126,
123, 127,
123, 128,
123, 165,
123, 166,
123, 167,
124, 125,
124, 126,
124, 127,
124, 128,
124, 129,
124, 167,
125, 126,
125, 127,
125, 128,
125, 129,
125, 130,
125, 132,
125, 147,
125, 150,
125, 151,
125, 154,
126, 127,
126, 128,
126, 129,
126, 130,
127, 128,
127, 129,
127, 130,
127, 131,
127, 132,
128, 129,
128, 130,
128, 131,
128, 132,
128, 147,
128, 150,
128, 154,
129, 143,
129, 147,
129, 150,
129, 151,
129, 130,
129, 131,
129, 132,
129, 133,
130, 131,
130, 132,
130, 133,
130, 134,
131, 132,
131, 133,
131, 134,
132, 133,
132, 134,
132, 143,
132, 146,
132, 147,
132, 150,
133, 143,
133, 146,
133, 147,
133, 134,
133, 135,
133, 136,
133, 137,
133, 138,
133, 140,
134, 143,
134, 135,
134, 136,
134, 137,
134, 138,
135, 136,
135, 137,
136, 143,
136, 137,
136, 138,
136, 139,
136, 140,
137, 138,
137, 139,
138, 141,
138, 142,
138, 143,
138, 146,
138, 139,
138, 140,
139, 140,
139, 141,
139, 142,
139, 143,
140, 141,
140, 142,
140, 143,
140, 144,
141, 142,
141, 143,
141, 144,
141, 145,
142, 143,
142, 144,
142, 145,
142, 146,
142, 147,
143, 144,
143, 145,
143, 146,
143, 147,
144, 145,
144, 146,
144, 147,
144, 148,
145, 146,
145, 147,
145, 148,
145, 149,
146, 147,
146, 148,
146, 149,
146, 150,
147, 148,
147, 149,
147, 150,
147, 151,
148, 149,
148, 150,
148, 151,
148, 152,
148, 153,
149, 150,
149, 151,
149, 152,
149, 153,
149, 154,
150, 151,
150, 152,
150, 153,
150, 154,
150, 155,
151, 152,
151, 153,
151, 154,
151, 155,
152, 153,
152, 154,
152, 155,
152, 156,
153, 154,
153, 155,
153, 156,
154, 155,
154, 156,
154, 157,
155, 156,
155, 157,
155, 158,
155, 159,
156, 157,
156, 158,
156, 159,
156, 160,
157, 158,
157, 159,
157, 160,
157, 163,
158, 159,
158, 160,
158, 161,
158, 163,
159, 160,
159, 161,
160, 161,
160, 162,
160, 163,
161, 162,
161, 163,
162, 163,
162, 164,
162, 179,
163, 164,
163, 165,
163, 175,
164, 165,
164, 166,
164, 167,
164, 172,
164, 175,
164, 176,
165, 166,
165, 167,
165, 171,
165, 172,
165, 175,
166, 167,
166, 168,
166, 169,
166, 171,
166, 172,
167, 168,
167, 171,
167, 172,
168, 169,
168, 170,
168, 171,
168, 172,
169, 170,
169, 171,
169, 172,
169, 173,
169, 174,
170, 171,
170, 172,
170, 173,
170, 174,
171, 172,
171, 173,
171, 174,
171, 175,
171, 176,
172, 173,
172, 174,
172, 175,
172, 176,
172, 177,
173, 174,
173, 175,
173, 176,
173, 177,
173, 178,
174, 175,
174, 176,
174, 177,
174, 178,
174, 182,
175, 176,
175, 177,
175, 178,
175, 179,
176, 177,
176, 178,
176, 179,
176, 180,
177, 178,
177, 179,
177, 180,
177, 181,
177, 182,
178, 179,
178, 180,
178, 181,
178, 182,
179, 180,
179, 181,
179, 182,
180, 181,
180, 182,
181, 182;
	springsstiffness = 
25.08,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01,
25.01;
	springsequilibrium = 
4.34437,
5.95684,
7.23055,
5.83643,
8.67239,
8.29299,
5.27912,
6.5669,
5.912,
4.95622,
6.07186,
7.68556,
8.79751,
6.58455,
4.69554,
7.52699,
7.98797,
4.85832,
5.585,
5.19389,
6.25207,
5.56837,
6.75822,
7.70859,
6.58126,
8.75401,
5.41901,
5.3163,
7.51841,
7.35018,
7.56628,
7.39957,
6.91409,
4.59699,
6.44124,
8.8232,
7.05713,
7.18101,
4.83872,
5.62043,
8.77459,
8.9863,
7.86169,
7.20221,
8.85903,
7.76626,
7.678,
4.48493,
5.0552,
5.77036,
4.41443,
5.93151,
7.29639,
5.27215,
7.19097,
6.17366,
7.40136,
7.06377,
6.25057,
8.64861,
5.81775,
7.18713,
4.7439,
8.14629,
6.48882,
5.09258,
7.99921,
6.56228,
5.815,
6.61228,
8.34676,
6.77899,
5.65806,
4.83325,
5.62704,
8.18603,
8.81593,
8.54118,
6.74294,
6.56406,
5.8885,
6.62273,
4.00106,
8.94439,
7.32073,
5.70232,
8.82876,
7.73728,
7.05642,
7.71035,
4.86019,
8.02943,
6.64498,
8.0629,
7.39865,
6.04187,
7.14634,
6.23594,
7.52694,
3.6655,
6.88158,
8.33666,
5.84921,
7.45044,
5.52466,
5.30911,
5.78343,
8.87016,
7.1189,
8.09492,
7.30356,
5.77133,
3.31354,
6.09949,
8.25585,
6.2721,
8.51418,
6.38119,
8.40983,
5.0465,
5.78383,
7.52213,
5.76545,
7.83878,
8.25842,
8.41714,
7.95948,
3.99054,
6.11794,
4.84673,
8.17871,
7.74741,
6.658,
6.70511,
6.9314,
7.3466,
7.67833,
8.68417,
6.29848,
4.55055,
6.18698,
3.75391,
5.64374,
7.9933,
7.84145,
7.54937,
7.75684,
8.01541,
7.87106,
6.73042,
6.19609,
4.24362,
5.7397,
7.68872,
6.3649,
6.34627,
6.88397,
3.92591,
6.18683,
8.60647,
8.82083,
8.61481,
5.25566,
6.01132,
6.05042,
8.77204,
6.93486,
8.13067,
6.43996,
4.73278,
5.1306,
4.91605,
5.99391,
8.29123,
6.45634,
8.66091,
6.5689,
7.78065,
5.4607,
7.81591,
4.55661,
7.09941,
6.54209,
6.38613,
6.51414,
6.97515,
3.74992,
5.43671,
4.69139,
6.47244,
8.49833,
4.44086,
6.20474,
5.67113,
6.81926,
8.95475,
6.01442,
4.43486,
7.3162,
5.29225,
5.84832,
7.65972,
7.87316,
5.85246,
8.74496,
6.58986,
5.59559,
7.57395,
6.44289,
6.3184,
6.16844,
6.07895,
5.33371,
6.2714,
8.7966,
7.41078,
8.65021,
5.30812,
8.01949,
6.78702,
5.52893,
4.10999,
7.34906,
4.71914,
4.98779,
8.23417,
7.14043,
7.91241,
8.73079,
5.47985,
8.60269,
8.92565,
6.9781,
6.44651,
6.93123,
6.17384,
5.87699,
7.17456,
8.85889,
5.56059,
8.02948,
6.419,
6.42616,
7.53522,
7.31857,
6.22161,
7.36244,
7.62705,
5.92413,
8.80722,
5.64767,
5.34209,
7.70737,
7.76035,
6.47019,
8.58066,
8.73795,
6.64771,
7.58852,
7.36765,
7.12748,
4.54155,
5.68579,
4.80804,
6.96453,
7.32775,
7.36555,
4.84245,
6.30129,
4.8487,
8.07734,
8.56367,
5.78442,
5.58672,
6.07289,
5.57987,
6.81269,
7.57537,
7.19587,
4.80674,
6.02083,
6.74756,
8.09772,
5.61267,
5.37954,
7.63572,
6.51362,
6.31683,
8.29982,
6.20334,
8.93886,
7.03105,
6.67297,
4.84786,
4.90982,
6.41389,
7.15029,
3.78246,
5.25707,
8.31097,
7.57415,
6.37019,
5.21453,
7.80612,
4.0076,
6.03559,
8.96071,
8.70106,
8.53577,
6.42371,
7.64542,
7.28775,
7.341,
7.34042,
8.88608,
3.91635,
6.92381,
5.65684,
6.82223,
7.22447,
6.13138,
5.64651,
8.23665,
7.93303,
7.94481,
8.47733,
3.45687,
6.4181,
7.55781,
8.2469,
4.59867,
5.22609,
8.51055,
6.63469,
4.73906,
6.08161,
6.67303,
4.07536,
7.38297,
8.81691,
8.75544,
5.68245,
4.94095,
7.24817,
6.41773,
6.63523,
8.35449,
5.14539,
4.01507,
6.74452,
6.14825,
5.38058,
6.99396,
5.33885,
5.69382,
8.57291,
7.18798,
8.86472,
6.61854,
7.87783,
5.49447,
6.9816,
4.17064,
5.00332,
7.45259,
8.87927,
7.69075,
5.80049,
6.46528,
4.96904,
6.36471,
8.78071,
8.51701,
5.42657,
5.87081,
7.05346,
5.95039,
7.21521,
6.68615,
6.06356,
8.96294,
5.98183,
8.98754,
3.81658,
5.62566,
6.24859,
8.07306,
6.12566,
8.72727,
3.4192,
7.03501,
8.12626,
8.96186,
5.5688,
5.90881,
6.67813,
7.41208,
5.29073,
8.5139,
8.73007,
8.34962,
8.58674,
5.71213,
7.62506,
5.12076,
4.62923,
6.04502,
8.28624,
4.25663,
6.12806,
7.88459,
4.98464,
7.46479,
7.07485,
5.18911,
7.98634,
4.93375,
5.93407,
4.7439,
5.26502,
8.9122,
7.6552,
6.33711,
7.21134,
8.20294,
5.60738,
5.06438,
8.97653,
4.14645,
3.66649,
5.74565,
6.99596,
4.48598,
7.21816,
4.11822,
7.73243,
7.84437,
4.89209,
8.16779,
7.50725,
6.28632,
5.93133,
8.04508,
8.23422,
5.97109,
6.86181,
8.37274,
6.90161,
8.80662,
6.1324,
5.02823,
6.53406,
8.58223,
6.26041,
6.19714,
8.83857,
3.44372,
4.94321,
6.46433,
7.58531,
8.79829,
4.38396,
7.97783,
6.30135,
7.6139,
8.8632,
7.14381,
6.35142,
7.41854,
5.89967,
5.4361,
8.88113,
6.7143,
8.08667,
4.81073,
4.99441,
8.38241,
5.7585,
7.686,
5.72403,
6.0604,
6.68903,
7.21494,
8.77375,
5.58599,
6.72712,
6.99531,
8.51186,
5.21764,
6.72404,
4.62305,
5.45595,
8.71362,
8.50723,
7.6609,
5.25956,
7.2492,
6.1731,
6.28155,
5.28738,
6.80041,
5.00136,
6.27138,
4.88715,
5.66311,
7.62518,
8.96821,
8.76482,
4.49303,
6.8999,
6.18653,
7.62353,
5.26797,
6.30818,
8.75092,
5.22682,
6.91396,
8.83156,
8.97644,
4.98071,
5.22002,
8.44948,
7.70051,
3.64189,
5.454,
7.24937,
7.47875,
5.40274,
7.61586,
6.71455,
5.28606,
5.8002,
8.66638,
5.11625,
5.9041,
6.7965,
8.7185,
6.20023,
5.66605,
5.52685,
6.56109,
8.1644,
6.39941,
4.70004,
8.99811,
4.84864,
6.86479,
5.12868,
8.05361,
4.94429,
6.94536,
5.53183,
8.01596,
7.51092,
8.49955,
7.72945,
5.20223,
7.68265,
6.13926,
6.21299,
8.83382,
5.99746,
6.86095,
7.35483,
5.183,
4.40875,
8.31721,
4.12905,
6.40993,
6.04612,
6.45905,
7.04225,
8.99408,
4.33899,
5.67624,
8.63387,
8.10232,
5.71452,
4.4811,
6.69244,
5.00211,
8.42676,
5.9043,
4.71213,
8.23124,
6.84123,
4.64417,
7.17216,
4.52787,
6.12146,
5.77923,
6.70038,
4.11499,
6.81254,
6.11057,
5.59584,
6.60233,
5.57011,
5.76321,
3.37012,
5.84849,
7.64854,
4.2486,
5.7307,
6.5352,
4.60517,
8.55578,
6.04018,
6.64111,
5.68305,
8.47713,
3.811,
7.72605,
4.00746,
6.04241,
7.26706,
8.48981,
8.46526,
7.3789,
4.62193,
6.63034,
8.44965,
8.19053,
4.60606,
5.91112,
5.68746,
7.58585,
8.3854,
8.38379,
4.33624,
5.20101,
5.08792,
5.96224,
8.38858,
4.79026,
7.26037,
7.59093,
7.3763,
4.36201,
7.67866,
5.76338,
6.85425,
8.25434,
7.68169,
5.06256,
5.83644,
5.52456,
6.43461,
8.84871,
6.29525,
6.3329,
7.82436,
6.06282,
7.21737,
5.9913,
7.12784,
7.70534,
3.50612,
5.19804,
4.94444,
5.62465,
8.23105,
3.53071,
5.11078,
4.73921,
5.67041,
4.48016,
6.8633,
6.65612,
3.58703,
5.3655,
5.09844,
5.84459,
7.65193,
7.42144,
7.34648,
3.82056,
5.65678,
5.15114,
8.85835,
4.08663,
3.44579,
6.1396,
8.92349,
3.85085,
6.75439,
7.86186,
5.87164,
7.11672,
4.64145,
4.9815,
6.41565,
7.1668,
4.51993,
7.04416,
7.71981,
5.93234,
6.17844,
8.45956,
7.6527,
4.84919,
8.50099,
4.40513,
7.09172,
7.23766,
5.26005,
5.87765,
8.19291,
4.30482,
4.38964,
4.85278,
6.29605,
8.81498,
4.8081,
6.36249,
5.89809,
6.9329,
7.89598,
6.47239,
6.76941,
7.36317,
3.37149,
5.04378,
5.44945,
6.20295,
8.43861,
3.22653,
6.45649,
4.63402,
5.52549,
5.36066,
5.11308,
4.85636,
6.88472,
8.65684,
6.4047,
7.44259,
5.65507,
8.15973,
8.93738,
7.22989,
6.70223,
6.9378,
8.03705,
8.91147,
4.09842,
6.67132,
4.77778,
6.04027,
8.96107,
5.75726,
7.10758,
5.47039,
6.03449,
8.03455,
7.20312,
8.38267,
5.83184,
7.06892,
6.41179,
4.5221,
7.4456,
5.38736,
7.5154,
6.60505,
7.78534,
5.5876,
8.89239,
7.49174,
5.03924,
6.5323,
8.61059,
4.53097,
4.1597,
5.06776,
8.99583,
4.11686,
5.4276,
8.98055,
4.51285,
8.16592,
7.71885,
4.04629,
6.5108,
4.32715,
6.1728,
8.40042,
5.32329,
6.60146,
7.49895,
4.60036,
8.02943,
7.84757,
4.33488,
4.24057,
6.6436,
8.9029,
5.96531,
6.836,
5.99604,
6.84769,
5.8115,
6.33175,
6.76808,
7.47611,
8.44158,
5.15745,
5.64138,
8.49722,
8.41062,
7.32559,
8.6565,
6.38947,
5.0794,
8.13983,
5.34034,
8.81017,
5.49512,
6.95781,
8.94197,
4.0966,
6.92831,
7.28783,
5.08742,
6.78521,
5.95191,
8.11645,
3.47666,
6.48553,
7.99475,
7.79562,
7.88915,
6.91862,
5.67267,
4.66915,
5.69535,
8.03049,
4.02163,
4.76519,
7.92707,
7.08373,
6.22218,
7.57476,
8.80607,
6.25782,
6.23433,
7.66237,
3.64128,
8.79485,
5.79754,
7.81968,
6.35632,
6.21756,
5.02656,
6.04341,
5.87762,
5.02596,
6.49059,
8.51174,
8.31834,
6.14662,
7.49723,
5.4835,
4.69607,
8.40282,
8.86562,
7.09982,
7.15332,
5.73146,
7.65535,
5.5247,
7.83281,
5.64812,
6.74517,
4.86692,
6.90242,
5.56382,
4.91946,
8.78747,
5.55255,
6.15163,
4.70904,
5.5332,
8.0086,
7.36834,
8.91892,
8.87406,
5.91084,
8.97702,
8.9422,
4.54795,
7.59906,
6.16008,
6.2678,
4.79316,
5.76599,
4.74258,
5.65983,
5.5664,
7.83452,
7.39732,
5.16514,
6.76341,
6.50318,
5.37484,
6.18223,
8.25643,
5.56466,
8.45027,
7.96694,
3.77072,
8.06529,
5.96461,
8.61096,
7.81787,
8.52489,
8.33811,
4.59511,
5.25415,
7.19028,
8.24258,
6.17984,
7.14333,
7.67228,
3.49898,
5.8942,
7.61427,
8.06727,
5.0629,
7.31791,
8.15125,
5.32236,
5.39542,
7.49559,
4.2537,
6.52822,
4.16865,
5.48507,
5.10226,
6.29676,
4.5249,
5.62444,
4.59743,
6.12301,
4.14299,
6.48564,
6.16497,
7.0461,
4.57273,
6.86283,
5.40557,
5.61804,
8.92726,
5.21334,
7.97776,
5.36381,
6.17183,
7.42788,
7.86201,
4.83528,
6.53465,
5.71023,
8.34906,
6.77614,
6.40499,
6.37239,
8.59818,
6.98013,
8.19941,
5.63077,
6.61974,
5.796,
6.98542,
4.11558,
5.9409,
6.72806,
5.8102,
8.63468,
4.10096,
8.104,
4.97693,
5.44811,
8.89798,
5.58957,
5.47539,
4.36094,
5.54355,
8.61534,
6.76712,
8.6331,
6.23336,
8.11018,
5.04275,
6.83404,
6.12596,
8.19239,
5.32849,
7.03238,
7.28252,
4.86074,
6.54106,
6.05429,
3.77226,
5.54768,
7.22033,
8.69386,
4.6061,
5.32052,
5.63718,
5.76536,
4.67442,
7.72373,
6.57389,
6.55572,
4.31149,
5.92692,
8.15088,
8.427,
4.82391,
7.187,
5.42546,
7.42586,
7.35742,
4.57935,
8.18315,
5.22701,
7.75554,
7.53187,
4.4264,
6.91034,
8.90977,
4.42143,
6.86069,
8.66617,
6.14994,
5.90022,
7.0345,
5.20248,
4.58584,
8.82844,
7.14682,
8.10816,
5.88922,
7.53143,
6.28587,
7.80718,
6.00106,
7.96471,
8.46191,
8.49635,
5.23536,
4.46151,
6.01915,
7.8414,
3.85423,
6.12795,
5.80104,
6.11395,
8.91177,
4.97484,
6.74337,
6.38398,
7.83372,
3.53434,
5.1717,
4.86482,
6.1992,
8.7308,
3.86517,
5.11297,
4.91484,
6.11585,
8.60157,
3.76147,
6.56224,
5.37805,
6.07697,
8.85745,
4.91496,
5.87813,
4.75655,
6.41593,
8.94854,
5.15925,
7.26648,
6.37933,
7.5945,
5.09421,
6.06741,
5.36187,
6.08889,
4.13885,
6.5716,
5.30015,
5.52225,
5.9394,
4.51885,
6.06371,
5.67339,
3.63958,
4.61255,
7.06736,
6.9095,
4.68999,
7.21312,
4.17768;
}
