netcdf SpringNetwork {

dimensions:
	spatialdim = 3;
	particle_number = 172;
	particlename_length = 5;
	chainname_length = 4;
	resname_length = 4;

variables:
	float   coordinates(particle_number, spatialdim); 
	        coordinates:units = "angstrom" ;
	        coordinates:long_name = "Particle coordinates";

	int     particleids(particle_number); 
	        particleids:long_name = "Particle ids in source database";

	char    particlenames(particle_number,particlename_length); 
	        particlenames:long_name = "Particle name";

	float   charges(particle_number);
	        charges:long_name = "Particle charge id";
	        charges:units = "electron" ;

	float   radii(particle_number);
	        radii:units = "A" ;
	        radii:long_name = "Particle radius";

	float   epsilon(particle_number);
	        epsilon:units = "kJ.mol-1" ;
	        epsilon:long_name = "Particle epsilon for Lennard-Jones";

	float   mass(particle_number);
	        mass:units = "Da" ;
	        mass:long_name = "Particle mass";

	float   surfaceaccessibility(particle_number);
	        surfaceaccessibility:units = "A2 or percent" ;
	        surfaceaccessibility:long_name = "Particle surface accessibility";

	float   hydrophobicityscale(particle_number);
	        hydrophobicityscale:units = "kJ.mol-1" ;
	        hydrophobicityscale:long_name = "Particle hydrophobicity scale (transfer energy)";

	char    resnames(particle_number,resname_length); 
	        resnames:long_name = "particle residue name";

	int     resids(particle_number); 
	        resids:long_name = "particle residue id";

	char    chainnames(particle_number,chainname_length); 
	        chainnames:long_name = "Chain name ";

	byte    dynamicstate(particle_number); 
	        dynamicstate:long_name = "particle dynamic state (static 0 or dynamic 1)";

	int     nbspringsperparticle(particle_number); 
	        nbspringsperparticle:long_name = "Number of springs per particle";

data:
	particleids = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	coordinates = 
-2.66812, -3.92325, -18.8477,
0.8478, -3.668, -16.7856,
2.25129, -0.833429, -16.2137,
3.34389, 0.750889, -21.1579,
8.24988, -1.62775, -20.007,
10.5778, 2.1155, -18.7859,
6.318, 3.72129, -17.133,
7.6135, 6.75507, -13.1459,
2.75217, 3.33417, -10.8632,
0.104571, 7.67029, -9.27371,
-2.1405, 6.6025, -6.135,
-5.002, 6.118, -4.0056,
-4.77078, 3.20533, -0.318889,
-9.66237, 4.15625, 0.8715,
-8.63675, 1.71725, 4.50025,
-11.0901, -2.287, 5.09479,
-7.97383, -2.348, 10.1763,
-11.3297, -5.21933, 12.3863,
-7.52592, -6.8765, 14.8455,
-3.182, -2.745, 12.9278,
-3.90112, -3.02975, 18.407,
-5.05829, -4.961, 21.409,
-4.511, -3.99425, 25.459,
-6.56812, -5.5575, 28.0389,
-6.69812, -4.0215, 32.9183,
-7.76937, -8.19312, 34.7181,
-10.312, -5.67912, 34.6784,
-12.3923, -5.58875, 30.2821,
-12.1308, -1.26825, 28.5217,
-12.0611, -1.43843, 25.2703,
-15.6851, -3.283, 23.0981,
-14.2333, -5.3483, 19.9191,
-10.0717, -1.79189, 17.5074,
-12.7662, -0.397, 13.789,
-7.98478, 0.881444, 12.7506,
-10.8269, 3.71088, 8.73687,
-7.8645, 5.03425, 5.8,
-5.446, 6.536, 3.6934,
-3.1925, 6.6445, 0.7395,
-0.312, 7.2724, -1.3762,
0.0964545, 4.25973, -4.82018,
4.28325, 5.22375, -6.3335,
5.8355, 4.0845, -9.51525,
10.0011, 2.55758, -13.0951,
6.55622, -1.14078, -14.1268,
10.959, -2.53086, -15.1513,
9.12925, -5.756, -16.4906,
5.61329, -7.00586, -17.4509,
6.32592, -10.2273, -15.5909,
9.05586, -5.98657, -12.1977,
8.136, -3.09625, -9.694,
10.6565, -1.325, -7.97655,
5.26833, 0.692333, -5.20833,
7.24662, 5.1545, -2.35588,
4.27675, 4.7945, 0.26925,
1.67658, 8.4055, 3.88975,
-0.149625, 4.35212, 4.53387,
-3.99371, 8.63829, 6.23271,
-4.5935, 3.89475, 9.97087,
-7.54625, 5.614, 12.4683,
-8.77218, 4.02018, 17.6104,
-13.1923, 5.31, 14.209,
-15.0506, 6.67157, 17.196,
-18.9755, 3.57692, 18.6356,
-19.1466, 2.25967, 23.1094,
-18.1012, 2.73675, 26.4853,
-16.744, 1.98683, 29.5703,
-14.8493, 4.75386, 31.5713,
-12.1479, 4.48867, 30.6963,
-10.0224, 4.56638, 25.2367,
-8.57125, 7.118, 22.8288,
-6.3708, 8.5384, 20.4148,
-3.7335, 4.4425, 17.1017,
-2.65422, 8.76811, 13.7946,
-0.8662, 5.4866, 12.1506,
1.86989, 8.03878, 9.961,
3.728, 5.3, 6.7025,
6.97143, 5.38214, 4.70957,
5.48167, 1.41656, 1.86556,
10.4605, 0.8225, -0.579,
7.84, -2.15186, -2.28857,
8.732, -4.8926, -4.672,
4.753, -4.73644, -8.14044,
6.55925, -9.38475, -8,
3.56275, -10.0443, -11.3577,
1.1635, -14.1524, -14.2607,
-0.348429, -11.7539, -16.3656,
-4.4175, -13.8846, -14.8911,
-6.09329, -11.435, -17.9884,
-5.14638, -8.86887, -21.3841,
-7.701, -6.47388, -18.274,
-6.68213, -9.276, -13.8953,
-2.4195, -8.16988, -12.8575,
-2.01662, -11.7358, -9.5215,
-0.42425, -7.24492, -6.442,
3.20014, -9.68171, -4.379,
3.29991, -4.68264, -2.07564,
8.47475, -7.72075, -1.23487,
9.46025, -4.7725, 2.15075,
9.6155, -1.58325, 3.765,
6.89388, 0.477625, 6.7695,
9.267, 3.80114, 8.33314,
6.24221, 1.9185, 12.9079,
4.98591, 8.41545, 14.8714,
2.4588, 5.5716, 16.649,
0.964375, 9.08725, 17.662,
-1.00743, 7.305, 21.5979,
-4.27525, 11.359, 24.5922,
-4.17467, 9.037, 27.7558,
-7.044, 10.2708, 30.162,
-3.83143, 9.296, 32.8357,
-0.557, 7.42358, 31.8035,
-1.05675, 11.1462, 27.5947,
1.05133, 13.4023, 24.1359,
3.39175, 8.06525, 23.7652,
6.3816, 8.6233, 20.4602,
6.30425, 3.87862, 18.9476,
9.17857, 4.328, 16.132,
9.68525, 1.772, 13.2325,
11.6129, -0.522571, 10.9377,
8.74817, -3.29133, 9.33183,
8.844, -6.13014, 7.55386,
5.88071, -4.80057, 4.098,
5.14609, -8.88727, 3.54282,
1.2146, -7.678, -0.2358,
-1.81175, -8.8795, -1.7695,
-3.35275, -8.6145, -5.0915,
-6.04443, -7.72271, -7.77,
-3.86522, -3.93833, -10.6518,
-9.87358, -4.56858, -13.9996,
-7.4384, -2.4472, -16.264,
-10.7071, 0.043125, -16.2131,
-8.41286, 2.127, -18.9403,
-5.15086, 2.11, -20.6369,
-5.00578, 5.556, -18.7934,
-7.6645, 3.83912, -14.7674,
-6.3054, 1.0844, -12.194,
-8.63514, -0.883, -9.844,
-4.03491, -1.54436, -6.354,
-8.343, -5.66263, -3.79925,
-3.71378, -4.43689, -1.32111,
-4.07308, -8.38258, 3.58008,
-0.622, -4.06067, 3.74556,
1.11286, -9.4405, 5.16379,
3.27386, -6.25186, 9.183,
6.1445, -9.74375, 10.1164,
5.67163, -7.61775, 14.1266,
9.80262, -9.8225, 15.5991,
11.1505, -6.3975, 17.5005,
14.2171, -4.58887, 18.5781,
12.8618, -3.6758, 23.0452,
11.0001, -4.0997, 26.3127,
11.0683, -5.111, 27.4646,
11.002, -9.38638, 25.945,
8.81775, -9.44925, 22.5472,
5.18114, -10.032, 21.8829,
4.954, -8.67673, 19.6532,
0.414143, -8.04786, 17.3407,
0.70175, -5.61775, 12.6744,
-3.43625, -7.31563, 11.6186,
-4.2, -6.15525, 8.55975,
-4.44413, -2.64925, 5.42413,
-8.29925, -4.77838, 3.3165,
-7.14667, -1.836, 0.245167,
-10.2802, -0.287, -2.23487,
-7.664, 1.4595, -5.4475,
-7.34571, 4.32286, -7.99457,
-4.01133, 4.04233, -10.6098,
-2.99225, 8.40483, -14.5239,
-1.37664, 2.88591, -15.7239,
1.81564, 9.16909, -15.5992,
2.95375, 6.46025, -20.205;
	charges = 
0,
0,
0,
1,
-1,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
1,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
-1,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
-1,
0,
0,
0,
1,
0,
0,
0,
1,
0,
0,
0,
-1,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
-1,
-1,
0,
-1,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
1,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
1,
0,
1,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
1,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
1,
0,
0,
0,
0,
1,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0;
	radii = 
3.47,
2.88,
3.2,
3.44,
3,
3.13,
3.12,
3.85,
3.66,
3.12,
2.58,
2.88,
3.44,
3.49,
2.58,
3.85,
2.89,
3.34,
3.66,
3.38,
3,
3.12,
2.58,
3.49,
3.47,
3.13,
3.13,
3.13,
2.58,
3.2,
3.12,
3.38,
3.22,
3.13,
3.44,
3.49,
2.58,
2.88,
2.58,
2.88,
3.64,
2.58,
2.58,
3.66,
3.34,
3.3,
3.13,
3.2,
3.66,
3.3,
2.58,
3.64,
3.22,
3.47,
2.58,
3.66,
3,
3.85,
3.49,
2.58,
3.47,
3.47,
3.2,
3.66,
3.44,
2.58,
2.89,
3.3,
3.22,
3.13,
2.58,
2.88,
3.66,
3.44,
2.88,
3.34,
2.58,
3.3,
3.34,
3.49,
3.12,
2.88,
3.44,
3.49,
2.58,
3.66,
3.2,
3.47,
3.12,
3,
3,
3.49,
3,
3.47,
3.66,
3.12,
3.47,
3.49,
2.58,
2.58,
3.47,
3.3,
3.85,
3.47,
2.88,
3,
3.12,
3.66,
2.89,
3.13,
3.3,
3.66,
2.58,
3.44,
3.13,
3.38,
3,
3.12,
2.58,
3.3,
2.89,
3.2,
3.3,
3.64,
2.88,
2.58,
2.58,
3.3,
3.22,
3.66,
2.88,
3.47,
3.12,
3.2,
3.22,
3.47,
2.88,
3.12,
3.47,
3.49,
3.22,
3.66,
3.34,
3.85,
3.12,
3.13,
3.13,
3.47,
2.58,
3,
2.88,
3.38,
3.12,
3.47,
2.58,
3.12,
3.47,
3.2,
3,
3.13,
2.58,
3.47,
3.49,
2.89,
3.49,
2.58,
3.3,
2.89,
3.66,
3.47,
3.64,
2.58;
	epsilon = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	mass = 
149,
89,
115,
146,
133,
132,
119,
204,
181,
119,
75,
89,
146,
131,
75,
204,
105,
146,
181,
155,
133,
119,
75,
131,
131,
132,
132,
132,
75,
115,
119,
155,
147,
132,
146,
131,
75,
89,
75,
89,
165,
75,
75,
181,
146,
117,
132,
115,
181,
117,
75,
165,
147,
149,
75,
181,
133,
204,
131,
75,
174,
149,
115,
181,
146,
75,
105,
117,
147,
132,
75,
89,
181,
146,
89,
146,
75,
117,
146,
131,
119,
89,
146,
131,
75,
181,
115,
131,
119,
133,
133,
131,
133,
131,
181,
119,
174,
131,
75,
75,
149,
117,
204,
174,
89,
133,
119,
181,
105,
132,
117,
181,
75,
146,
132,
155,
133,
119,
75,
117,
105,
115,
117,
165,
89,
75,
75,
117,
147,
181,
89,
131,
119,
115,
147,
131,
89,
119,
174,
131,
147,
181,
146,
204,
119,
132,
132,
131,
75,
133,
89,
155,
119,
131,
75,
119,
174,
115,
133,
132,
75,
149,
131,
105,
131,
75,
117,
105,
181,
174,
165,
75;
	surfaceaccessibility = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	hydrophobicityscale = 
0.026388,
0.011407,
0.021775,
-0.020395,
-0.022949,
-0.017252,
0.007727,
0.036833,
0.018661,
0.007727,
0,
0.011407,
-0.020395,
0.038397,
0,
0.036833,
-0.001417,
-0.005096,
0.018661,
0.002943,
-0.022949,
0.007727,
0,
0.038397,
0.042811,
-0.017252,
-0.017252,
-0.017252,
0,
0.021775,
0.007727,
0.002943,
-0.015356,
-0.017252,
-0.020395,
0.038397,
0,
0.011407,
0,
0.011407,
0.037028,
0,
0,
0.018661,
-0.005096,
0.033514,
-0.017252,
0.021775,
0.018661,
0.033514,
0,
0.037028,
-0.015356,
0.026388,
0,
0.018661,
-0.022949,
0.036833,
0.038397,
0,
-0.017504,
0.026388,
0.021775,
0.018661,
-0.020395,
0,
-0.001417,
0.033514,
-0.015356,
-0.017252,
0,
0.011407,
0.018661,
-0.020395,
0.011407,
-0.005096,
0,
0.033514,
-0.005096,
0.038397,
0.007727,
0.011407,
-0.020395,
0.038397,
0,
0.018661,
0.021775,
0.042811,
0.007727,
-0.022949,
-0.022949,
0.038397,
-0.022949,
0.042811,
0.018661,
0.007727,
-0.017504,
0.038397,
0,
0,
0.026388,
0.033514,
0.036833,
-0.017504,
0.011407,
-0.022949,
0.007727,
0.018661,
-0.001417,
-0.017252,
0.033514,
0.018661,
0,
-0.020395,
-0.017252,
0.002943,
-0.022949,
0.007727,
0,
0.033514,
-0.001417,
0.021775,
0.033514,
0.037028,
0.011407,
0,
0,
0.033514,
-0.015356,
0.018661,
0.011407,
0.042811,
0.007727,
0.021775,
-0.015356,
0.042811,
0.011407,
0.007727,
-0.017504,
0.038397,
-0.015356,
0.018661,
-0.005096,
0.036833,
0.007727,
-0.017252,
-0.017252,
0.042811,
0,
-0.022949,
0.011407,
0.002943,
0.007727,
0.042811,
0,
0.007727,
-0.017504,
0.021775,
-0.022949,
-0.017252,
0,
0.026388,
0.038397,
-0.001417,
0.038397,
0,
0.033514,
-0.001417,
0.018661,
-0.017504,
0.037028,
0;
	particlenames = 
"MCA",
"ACA",
"PCA",
"KCA",
"DCA",
"NCA",
"TCA",
"WCA",
"YCA",
"TCA",
"GCA",
"ACA",
"KCA",
"LCA",
"GCA",
"WCA",
"SCA",
"QCA",
"YCA",
"HCA",
"DCA",
"TCA",
"GCA",
"LCA",
"ICA",
"NCA",
"NCA",
"NCA",
"GCA",
"PCA",
"TCA",
"HCA",
"ECA",
"NCA",
"KCA",
"LCA",
"GCA",
"ACA",
"GCA",
"ACA",
"FCA",
"GCA",
"GCA",
"YCA",
"QCA",
"VCA",
"NCA",
"PCA",
"YCA",
"VCA",
"GCA",
"FCA",
"ECA",
"MCA",
"GCA",
"YCA",
"DCA",
"WCA",
"LCA",
"GCA",
"RCA",
"MCA",
"PCA",
"YCA",
"KCA",
"GCA",
"SCA",
"VCA",
"ECA",
"NCA",
"GCA",
"ACA",
"YCA",
"KCA",
"ACA",
"QCA",
"GCA",
"VCA",
"QCA",
"LCA",
"TCA",
"ACA",
"KCA",
"LCA",
"GCA",
"YCA",
"PCA",
"ICA",
"TCA",
"DCA",
"DCA",
"LCA",
"DCA",
"ICA",
"YCA",
"TCA",
"RCA",
"LCA",
"GCA",
"GCA",
"MCA",
"VCA",
"WCA",
"RCA",
"ACA",
"DCA",
"TCA",
"YCA",
"SCA",
"NCA",
"VCA",
"YCA",
"GCA",
"KCA",
"NCA",
"HCA",
"DCA",
"TCA",
"GCA",
"VCA",
"SCA",
"PCA",
"VCA",
"FCA",
"ACA",
"GCA",
"GCA",
"VCA",
"ECA",
"YCA",
"ACA",
"ICA",
"TCA",
"PCA",
"ECA",
"ICA",
"ACA",
"TCA",
"RCA",
"LCA",
"ECA",
"YCA",
"QCA",
"WCA",
"TCA",
"NCA",
"NCA",
"ICA",
"GCA",
"DCA",
"ACA",
"HCA",
"TCA",
"ICA",
"GCA",
"TCA",
"RCA",
"PCA",
"DCA",
"NCA",
"GCA",
"MCA",
"LCA",
"SCA",
"LCA",
"GCA",
"VCA",
"SCA",
"YCA",
"RCA",
"FCA",
"GCA";
	resnames = 
"MET",
"ALA",
"PRO",
"LYS",
"ASP",
"ASN",
"THR",
"TRP",
"TYR",
"THR",
"GLY",
"ALA",
"LYS",
"LEU",
"GLY",
"TRP",
"SER",
"GLN",
"TYR",
"HIS",
"ASP",
"THR",
"GLY",
"LEU",
"ILE",
"ASN",
"ASN",
"ASN",
"GLY",
"PRO",
"THR",
"HIS",
"GLU",
"ASN",
"LYS",
"LEU",
"GLY",
"ALA",
"GLY",
"ALA",
"PHE",
"GLY",
"GLY",
"TYR",
"GLN",
"VAL",
"ASN",
"PRO",
"TYR",
"VAL",
"GLY",
"PHE",
"GLU",
"MET",
"GLY",
"TYR",
"ASP",
"TRP",
"LEU",
"GLY",
"ARG",
"MET",
"PRO",
"TYR",
"LYS",
"GLY",
"SER",
"VAL",
"GLU",
"ASN",
"GLY",
"ALA",
"TYR",
"LYS",
"ALA",
"GLN",
"GLY",
"VAL",
"GLN",
"LEU",
"THR",
"ALA",
"LYS",
"LEU",
"GLY",
"TYR",
"PRO",
"ILE",
"THR",
"ASP",
"ASP",
"LEU",
"ASP",
"ILE",
"TYR",
"THR",
"ARG",
"LEU",
"GLY",
"GLY",
"MET",
"VAL",
"TRP",
"ARG",
"ALA",
"ASP",
"THR",
"TYR",
"SER",
"ASN",
"VAL",
"TYR",
"GLY",
"LYS",
"ASN",
"HIS",
"ASP",
"THR",
"GLY",
"VAL",
"SER",
"PRO",
"VAL",
"PHE",
"ALA",
"GLY",
"GLY",
"VAL",
"GLU",
"TYR",
"ALA",
"ILE",
"THR",
"PRO",
"GLU",
"ILE",
"ALA",
"THR",
"ARG",
"LEU",
"GLU",
"TYR",
"GLN",
"TRP",
"THR",
"ASN",
"ASN",
"ILE",
"GLY",
"ASP",
"ALA",
"HIS",
"THR",
"ILE",
"GLY",
"THR",
"ARG",
"PRO",
"ASP",
"ASN",
"GLY",
"MET",
"LEU",
"SER",
"LEU",
"GLY",
"VAL",
"SER",
"TYR",
"ARG",
"PHE",
"GLY";
	resids = 
0,
1,
2,
3,
4,
5,
6,
7,
8,
9,
10,
11,
12,
13,
14,
15,
16,
17,
18,
19,
20,
21,
22,
23,
24,
25,
26,
27,
28,
29,
30,
31,
32,
33,
34,
35,
36,
37,
38,
39,
40,
41,
42,
43,
44,
45,
46,
47,
48,
49,
50,
51,
52,
53,
54,
55,
56,
57,
58,
59,
60,
61,
62,
63,
64,
65,
66,
67,
68,
69,
70,
71,
72,
73,
74,
75,
76,
77,
78,
79,
80,
81,
82,
83,
84,
85,
86,
87,
88,
89,
90,
91,
92,
93,
94,
95,
96,
97,
98,
99,
100,
101,
102,
103,
104,
105,
106,
107,
108,
109,
110,
111,
112,
113,
114,
115,
116,
117,
118,
119,
120,
121,
122,
123,
124,
125,
126,
127,
128,
129,
130,
131,
132,
133,
134,
135,
136,
137,
138,
139,
140,
141,
142,
143,
144,
145,
146,
147,
148,
149,
150,
151,
152,
153,
154,
155,
156,
157,
158,
159,
160,
161,
162,
163,
164,
165,
166,
167,
168,
169,
170,
171;
	chainnames = 
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A";
	dynamicstate = 
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1;
	nbspringsperparticle = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
}
