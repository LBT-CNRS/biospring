netcdf SpringNetwork {

dimensions:
	spatialdim = 3;
	particle_number = 397;
	particlename_length = 5;
	chainname_length = 4;
	resname_length = 4;

	springdim = 2; 
	spring_number = 1072;

variables:
	float   coordinates(particle_number, spatialdim); 
	        coordinates:units = "angstrom" ;
	        coordinates:long_name = "Particle coordinates";

	int     particleids(particle_number); 
	        particleids:long_name = "Particle ids in source database";

	char    particlenames(particle_number,particlename_length); 
	        particlenames:long_name = "Particle name";

	float   charges(particle_number);
	        charges:long_name = "Particle charge id";
	        charges:units = "electron" ;

	float   radii(particle_number);
	        radii:units = "A" ;
	        radii:long_name = "Particle radius";

	float   epsilon(particle_number);
	        epsilon:units = "kJ.mol-1" ;
	        epsilon:long_name = "Particle epsilon for Lennard-Jones";

	float   mass(particle_number);
	        mass:units = "Da" ;
	        mass:long_name = "Particle mass";

	float   surfaceaccessibility(particle_number);
	        surfaceaccessibility:units = "A2 or percent" ;
	        surfaceaccessibility:long_name = "Particle surface accessibility";

	float   hydrophobicityscale(particle_number);
	        hydrophobicityscale:units = "kJ.mol-1" ;
	        hydrophobicityscale:long_name = "Particle hydrophobicity scale (transfer energy)";

	char    resnames(particle_number,resname_length); 
	        resnames:long_name = "particle residue name";

	int     resids(particle_number); 
	        resids:long_name = "particle residue id";

	char    chainnames(particle_number,chainname_length); 
	        chainnames:long_name = "Chain name ";

	byte    dynamicstate(particle_number); 
	        dynamicstate:long_name = "particle dynamic state (static 0 or dynamic 1)";

	int     nbspringsperparticle(particle_number); 
	        nbspringsperparticle:long_name = "Number of springs per particle";

	int     springs(spring_number,springdim); 
	        springs:long_name = "Spring between particle referenced by 2 particle ids"; 

	float   springsstiffness(spring_number); 
	        springsstiffness:long_name = "Spring stiffness";
	float   springsequilibrium(spring_number); 
	        springsequilibrium:long_name = "Spring distance equilibrium";
data:
	particleids = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	coordinates = 
-2.069, -4.848, -17.494,
-3.268, -2.998, -20.201,
0.848, -3.668, -16.786,
2.506, -1.139, -17.159,
1.912, -0.426, -14.953,
4.668, 0.111, -19.197,
3.241, 0.952, -22.153,
0.849, 1.729, -23.587,
7.957, -0.294, -19.251,
8.543, -2.962, -20.763,
9.276, 2.942, -18.515,
11.879, 1.289, -19.057,
6.943, 3.696, -16.213,
5.485, 3.756, -18.36,
4.683, 5.596, -14.357,
6.671, 7.18, -13.551,
8.812, 7.537, -14.58,
8.988, 7.261, -12.799,
8.767, 6.898, -10.768,
10.691, 7.217, -11.609,
2.72, 5.835, -11.272,
1.865, 3.648, -11.807,
3.559, 1.883, -11.524,
1.986, 2.253, -9.742,
3.664, 0.551, -9.56,
-0.308, 6.663, -9.383,
0.654, 9.014, -9.128,
-2.14, 6.603, -6.135,
-5.002, 6.118, -4.006,
-6.402, 4.762, -0.829,
-4.334, 2.547, -0.635,
-2.163, 1.079, 1.175,
-8.621, 2.866, 1.172,
-10.704, 5.447, 0.571,
-8.637, 1.717, 4.5,
-8.975, -1.245, 6.664,
-11.335, -1.541, 6.375,
-11.848, -3.865, 6.014,
-11.985, -2.939, 4.474,
-12.036, -1.563, 2.919,
-12.476, -3.61, 2.554,
-8.774, -2.196, 10.135,
-6.374, -2.651, 10.259,
-9.863, -4.515, 12.666,
-12.503, -5.783, 12.162,
-7.027, -4.548, 14.194,
-7.982, -6.004, 15.792,
-6.587, -7.957, 15.217,
-8.963, -8.175, 15.118,
-7.571, -10.027, 14.558,
-3.628, -3.471, 15.02,
-3.38, -2.108, 12.913,
-1.946, -1.837, 11.023,
-3.329, -2.839, 10.663,
-4.067, -4.441, 18.024,
-3.735, -1.619, 18.79,
-4.118, -4.342, 21.769,
-6.312, -5.787, 20.929,
-4.511, -3.994, 25.459,
-5.546, -4.485, 28.897,
-7.59, -6.63, 27.181,
-7.112, -5.436, 32.312,
-6.284, -2.607, 33.524,
-7.849, -7.389, 33.198,
-7.69, -8.998, 36.238,
-10.067, -5.583, 33.094,
-10.557, -5.775, 36.263,
-11.914, -4.136, 30.88,
-12.87, -7.041, 29.684,
-12.131, -1.268, 28.522,
-12.927, -1.813, 25.495,
-10.907, -0.94, 24.971,
-14.754, -3.782, 22.902,
-16.927, -2.617, 23.36,
-13.378, -3.113, 20.048,
-14.588, -5.661, 19.492,
-14.094, -7.659, 19.72,
-15.728, -7.196, 20.286,
-11.893, -2.44, 16.615,
-8.614, -1.274, 18.222,
-11.42, 0.393, 14.28,
-14.113, -1.187, 13.297,
-9.69, 1.21, 11.239,
-7.28, 0.838, 13.136,
-5.631, 0.289, 15.196,
-9.209, 4.013, 9.102,
-12.445, 3.409, 8.372,
-7.865, 5.034, 5.8,
-5.446, 6.536, 3.693,
-3.193, 6.644, 0.74,
-0.312, 7.272, -1.376,
1.288, 6.037, -4.487,
0.462, 3.644, -4.215,
-1.813, 3.149, -4.796,
-0.643, 2.847, -6.204,
4.283, 5.224, -6.334,
5.835, 4.085, -9.515,
7.895, 1.768, -11.383,
9.86, 3.139, -12.191,
10.479, 3.87, -14.466,
11.653, 2.033, -13.477,
12.224, 2.767, -15.669,
8.154, 0.07, -14.309,
5.278, -2.11, -13.981,
10.131, -2.41, -15.881,
12.062, -2.692, -14.178,
8.14, -4.777, -16.501,
10.118, -6.735, -16.481,
5.387, -6.89, -16.436,
5.915, -7.16, -18.805,
6.49, -8.154, -13.491,
6.999, -10.211, -14.95,
5.393, -11.758, -15.971,
7.094, -10.778, -17.354,
5.49, -12.309, -18.289,
8.189, -5.405, -12.468,
10.212, -6.762, -11.838,
8.136, -3.096, -9.694,
8.381, -0.032, -7.812,
11.126, -1.037, -7.763,
12.314, -3.075, -7.434,
12.622, -2.316, -9.087,
7.245, 1.333, -4.574,
3.687, 0.18, -5.715,
5.798, 4.123, -2.983,
8.695, 6.186, -1.729,
4.277, 4.795, 0.269,
1.651, 6.314, 2.173,
2.434, 8.524, 2.982,
2.628, 9.043, 5.383,
0.74, 9.883, 4.155,
0.956, 10.355, 6.471,
0.027, 5.809, 5.333,
-0.326, 2.895, 3.735,
-3.101, 6.037, 7.228,
-3.089, 8.446, 7.328,
-5.349, 9.179, 7.418,
-4.574, 9.738, 5.88,
-3.377, 10.175, 4.246,
-5.367, 10.857, 4.3,
-4.505, 5.517, 10.559,
-4.682, 2.272, 9.383,
-7.546, 5.614, 12.468,
-9.361, 5.394, 15.104,
-9.257, 3.768, 17.647,
-7.82, 2.836, 20.089,
-12.693, 4.601, 15.748,
-13.691, 6.019, 12.67,
-15.346, 5.844, 17.492,
-14.657, 7.775, 16.802,
-16.443, 3.091, 19.871,
-18.287, 2.986, 18.185,
-20.613, 3.229, 18.998,
-19.915, 4.422, 17.049,
-22.151, 4.643, 17.838,
-16.59, 2.152, 22.917,
-19.962, 2.263, 23.429,
-23.038, 2.47, 23.016,
-18.101, 2.737, 26.485,
-16.707, 2.617, 29.828,
-16.819, 0.726, 29.055,
-14.721, 4.476, 30.576,
-15.021, 5.125, 32.899,
-11.803, 5.162, 28.717,
-12.424, 3.95, 32.28,
-10.846, 5.988, 25.163,
-9.199, 3.144, 25.311,
-8.571, 7.118, 22.829,
-6.371, 8.538, 20.415,
-5.239, 6.774, 17.223,
-4.51, 4.503, 17.923,
-3.433, 3.451, 15.946,
-2.493, 3.073, 18.117,
-1.486, 2.079, 16.178,
-2.332, 6.936, 15.094,
-2.826, 9.786, 13.801,
-3.041, 10.905, 11.186,
-0.866, 5.487, 12.151,
2.094, 5.857, 10.065,
1.69, 9.784, 9.878,
3.728, 5.3, 6.703,
6.59, 4.383, 4.851,
7.48, 6.715, 4.521,
7.164, 2.637, 1.766,
4.136, 0.44, 1.945,
9.245, 0.107, 0.047,
11.676, 1.538, -1.204,
8.71, -1.891, -2.931,
6.681, -2.5, -1.432,
8.732, -4.893, -4.672,
6.608, -5.724, -7.539,
3.861, -4.312, -7.765,
2.382, -3.397, -9.907,
4.994, -8.85, -8.245,
8.125, -9.919, -7.755,
3.563, -10.044, -11.358,
0.778, -11.677, -13.06,
1.637, -14.026, -13.255,
2.475, -15.184, -15.265,
0.236, -15.623, -14.491,
1.076, -16.728, -16.433,
-1.051, -12.128, -15.971,
0.588, -11.255, -16.891,
-4.162, -13.579, -16.16,
-4.673, -14.19, -13.622,
-4.978, -11.329, -18.187,
-7.58, -11.576, -17.724,
-5.129, -8.229, -19.916,
-5.164, -9.509, -22.853,
-6.578, -6.864, -17.187,
-8.823, -6.084, -19.361,
-5.486, -9.009, -14.874,
-7.879, -9.543, -12.916,
-3.627, -8.849, -11.896,
-1.212, -7.49, -13.819,
-1.389, -10.418, -9.757,
-2.645, -13.054, -9.285,
0.2, -9.62, -6.567,
0.51, -7.414, -7.474,
0.069, -6.005, -5.487,
-1.577, -6.082, -7.257,
-1.947, -4.729, -5.3,
3.111, -8.655, -4.796,
3.32, -11.05, -3.823,
4.657, -7.117, -2.009,
3.27, -4.299, -3.233,
1.966, -2.535, -1.274,
8.056, -6.313, -0.939,
8.893, -9.128, -1.531,
9.46, -4.772, 2.151,
9.615, -1.583, 3.765,
8.726, 0.206, 6.965,
5.061, 0.749, 6.574,
8.244, 3.361, 8.362,
10.631, 4.388, 8.294,
6.86, 4.041, 11.609,
5.601, 2.115, 11.406,
6.728, 0.065, 11.954,
6.111, 0.861, 13.447,
5.278, 2.065, 14.901,
6.258, 0.243, 15.43,
4.164, 5.807, 13.528,
5.37, 8.422, 14.31,
5.52, 11.019, 16.636,
2.459, 5.572, 16.649,
-0.001, 7.863, 18.165,
1.93, 10.312, 17.159,
-1.103, 8.43, 21.339,
-0.879, 5.805, 21.944,
-3.666, 8.572, 24.013,
-4.322, 11.071, 23.578,
-3.513, 13.175, 24.58,
-5.668, 12.361, 25.216,
-4.817, 14.402, 26.152,
-4.396, 9.765, 27.337,
-3.732, 7.58, 28.594,
-5.677, 10.975, 30.325,
-8.411, 9.567, 29.999,
-3.578, 10.271, 32.255,
-4.169, 7.995, 33.611,
-0.694, 10.037, 30.405,
-0.454, 7.553, 30.917,
0.377, 6.696, 33.083,
-1.364, 5.497, 31.957,
-0.513, 4.722, 34.053,
-1.057, 11.146, 27.595,
1.252, 11.428, 25.218,
0.487, 13.957, 23.265,
1.495, 16.52, 23.278,
2.457, 8.956, 22.795,
4.327, 7.175, 24.735,
5.055, 7.217, 21.022,
5.897, 9.127, 19.788,
8.203, 8.946, 20.382,
7.697, 10.61, 20.086,
6.246, 5.301, 18.163,
6.362, 2.456, 19.732,
8.742, 3.298, 16.487,
9.761, 5.701, 15.659,
9.685, 1.772, 13.232,
10.734, -1.106, 11.445,
12.785, 0.255, 10.261,
9.313, -3.068, 8.722,
7.619, -3.737, 10.552,
8.189, -5.55, 7.135,
9.718, -6.903, 8.113,
6.317, -5.806, 4.018,
5.3, -3.46, 4.204,
3.187, -7.205, 2.812,
5.03, -9.463, 3.507,
7.344, -10.069, 3.381,
6.707, -10.104, 5.097,
1.215, -7.678, -0.236,
-1.812, -8.88, -1.769,
-3.353, -8.614, -5.091,
-5.406, -6.84, -7.413,
-6.896, -8.9, -8.246,
-5.34, -5.54, -10.791,
-2.686, -2.657, -10.54,
-7.56, -3.474, -12.829,
-9.61, -4.916, -12.994,
-11.101, -3.948, -14.689,
-10.986, -6.316, -14.513,
-12.425, -5.285, -16.145,
-7.438, -2.447, -16.264,
-9.996, -0.411, -17.375,
-11.418, 0.497, -15.052,
-7.854, 1.212, -18.761,
-9.158, 3.347, -19.179,
-4.714, 2.194, -19.668,
-5.733, 1.997, -21.928,
-4.74, 4.555, -17.201,
-5.219, 6.357, -20.068,
-6.809, 2.9, -15.236,
-8.521, 4.778, -14.298,
-6.305, 1.084, -12.194,
-7.573, -1.118, -9.786,
-10.051, -0.57, -9.921,
-7.272, -2.207, -6.276,
-4.207, -1.536, -6.419,
-0.668, -0.889, -6.383,
-6.954, -5.134, -4.277,
-9.732, -6.191, -3.322,
-5.641, -5.293, -0.95,
-2.172, -3.752, -1.618,
-3.43, -6.985, 1.351,
-4.711, -8.627, 2.641,
-5.278, -8.338, 5.014,
-3.479, -9.851, 4.418,
-4.112, -9.509, 6.704,
-1.638, -5.889, 4.201,
0.191, -2.598, 3.381,
1.322, -6.858, 6.015,
0.417, -9.049, 6.544,
2.081, -10.774, 6.428,
1.203, -10.647, 4.857,
-0.007, -10.178, 3.209,
1.451, -11.721, 3.079,
3.072, -7.258, 9.056,
3.543, -4.91, 9.353,
5.52, -8.725, 10.793,
6.769, -10.762, 9.44,
5.548, -9.201, 14.581,
5.795, -6.034, 13.673,
9.066, -8.553, 16.318,
10.539, -11.091, 14.88,
11.151, -6.398, 17.5,
12.907, -4.045, 19.44,
15.527, -5.133, 17.716,
12.862, -3.676, 23.045,
12.44, -2.325, 26.432,
10.802, -4.182, 26.777,
9.01, -5.591, 26.509,
10.309, -6.077, 25.413,
12.037, -5.416, 26.977,
9.777, -4.704, 28.115,
10.104, -8.155, 25.486,
11.9, -10.617, 26.404,
8.818, -9.449, 22.547,
5.366, -9.656, 20.769,
4.935, -10.533, 23.368,
1.744, -9.14, 19.282,
4.963, -9.429, 18.876,
8.157, -7.649, 20.608,
0.476, -7.212, 17.159,
0.332, -9.162, 17.583,
0.303, -6.548, 13.636,
1.101, -4.688, 11.713,
-2.208, -6.312, 11.233,
-4.664, -8.319, 12.005,
-4.2, -6.155, 8.56,
-4.822, -4.385, 5.478,
-4.066, -0.913, 5.37,
-7.481, -3.34, 3.575,
-9.117, -6.216, 3.058,
-7.766, -2.255, 0.05,
-5.908, -0.998, 0.636,
-8.74, 0.328, -2.188,
-11.821, -0.902, -2.282,
-7.664, 1.46, -5.447,
-6.311, 3.99, -7.634,
-8.726, 4.767, -8.475,
-4.637, 4.471, -10.859,
-2.76, 3.186, -10.111,
-2.347, 6.33, -12.788,
-3.413, 8.469, -13.506,
-4.424, 9.069, -15.665,
-2.194, 9.83, -15.159,
-3.229, 10.401, -17.236,
-0.941, 6.176, -16.027,
-1.069, 2.987, -15.727,
-2.043, -0.48, -15.418,
2.013, 7.488, -17.549,
2.147, 9.516, -15.628,
1.127, 11.219, -14.28,
1.731, 9.797, -13.284,
3.029, 6.448, -20.608;
	charges = 
0,
0,
0,
0,
0,
0,
0,
1,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
-1,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
-1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
0,
0,
0,
0;
	radii = 
2.35,
2.35,
2.35,
2.05,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
1.7,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.35,
2.35,
2.05,
2.05,
2.35,
2.05,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
1.7,
2.35,
1.7,
2.35,
2.35,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
1.7,
1.7,
1.7,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.05,
2.05,
2.05,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
2.35,
2.35,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
2.35,
1.7,
1.7,
1.7,
2.05,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.35,
2.35,
2.05,
2.35,
2.05,
2.05,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.35,
1.7,
1.7,
1.7,
2.35,
2.35,
2.35,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.35,
2.05,
2.05,
2.35,
2.35,
2.05,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.05,
2.35,
1.7,
2.35,
2.05,
2.35,
2.35,
2.35,
2.05,
2.05,
2.35,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.35,
2.35,
2.35,
2.05,
2.35,
2.05,
2.35,
2.35,
2.35,
2.05,
2.35,
2.05,
2.35,
2.35,
2.05,
2.05,
2.35,
2.05,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.05,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.05,
2.05,
2.35,
2.35,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.35,
2.35,
2.05,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
1.7,
2.35,
2.05,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
1.7,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
1.7,
2.05,
2.05,
2.35,
2.05,
2.35,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
2.35,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.35,
2.05,
2.35,
2.05,
2.05,
2.05,
2.35,
2.35,
2.35,
2.05,
2.35,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
2.35,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.35,
2.35,
1.7,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
2.35,
1.7,
1.7,
1.7,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
2.05,
2.05,
2.05,
2.05,
2.35,
2.05,
2.35,
2.05,
2.05,
2.35,
2.35,
2.35,
2.05,
2.35,
1.7,
2.35,
2.05,
2.05,
2.35,
2.05,
2.35,
1.7,
2.35,
1.7,
1.7,
1.7,
1.7,
2.35,
2.05,
2.05,
2.35,
1.7,
1.7,
1.7,
2.05;
	epsilon = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	mass = 
72,
72,
72,
54,
54,
72,
54,
54,
72,
54,
72,
54,
72,
54,
72,
36,
36,
36,
36,
36,
72,
36,
36,
36,
36,
72,
54,
54,
72,
72,
54,
54,
72,
54,
54,
72,
36,
36,
36,
36,
36,
72,
36,
72,
72,
72,
36,
36,
36,
36,
72,
36,
36,
36,
72,
54,
72,
54,
54,
72,
54,
72,
54,
72,
54,
72,
54,
72,
54,
54,
54,
54,
72,
54,
72,
36,
36,
36,
72,
72,
72,
54,
72,
54,
54,
72,
54,
54,
72,
54,
72,
72,
36,
36,
36,
54,
54,
72,
36,
36,
36,
36,
72,
72,
72,
54,
72,
54,
54,
54,
72,
36,
36,
36,
36,
72,
54,
54,
72,
36,
36,
36,
72,
72,
72,
72,
54,
72,
36,
36,
36,
36,
72,
54,
72,
36,
36,
36,
36,
36,
72,
54,
54,
72,
54,
54,
72,
72,
54,
54,
72,
36,
36,
36,
36,
72,
54,
54,
54,
72,
36,
72,
54,
72,
72,
72,
54,
54,
72,
72,
36,
36,
36,
36,
72,
54,
54,
72,
72,
72,
54,
72,
54,
72,
72,
72,
54,
72,
54,
72,
72,
54,
54,
72,
54,
54,
72,
36,
36,
36,
36,
54,
54,
72,
54,
72,
54,
72,
54,
72,
54,
72,
54,
72,
54,
72,
54,
72,
36,
36,
36,
36,
72,
54,
72,
54,
54,
72,
54,
54,
54,
72,
72,
72,
54,
72,
36,
36,
36,
36,
36,
72,
54,
54,
72,
72,
54,
72,
54,
72,
36,
36,
36,
36,
72,
36,
72,
54,
72,
54,
72,
36,
36,
36,
36,
54,
72,
54,
54,
72,
54,
72,
36,
36,
36,
72,
54,
72,
54,
54,
72,
54,
72,
36,
54,
54,
72,
54,
72,
36,
36,
36,
72,
54,
54,
72,
54,
72,
72,
72,
36,
36,
36,
36,
72,
72,
54,
72,
54,
54,
54,
72,
72,
72,
54,
72,
72,
54,
72,
54,
54,
72,
54,
72,
72,
72,
36,
36,
36,
36,
72,
72,
72,
36,
36,
36,
36,
36,
72,
54,
72,
54,
72,
54,
72,
54,
54,
72,
54,
72,
72,
36,
36,
36,
72,
54,
72,
54,
54,
72,
54,
72,
54,
54,
54,
54,
72,
54,
72,
54,
54,
72,
72,
72,
54,
72,
36,
72,
54,
54,
72,
54,
72,
36,
72,
36,
36,
36,
36,
72,
54,
54,
72,
36,
36,
36,
54;
	surfaceaccessibility = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	hydrophobicityscale = 
0.0209,
-0.1029,
-0.065,
0.0307,
-0.0772,
0.0085,
-0.0337,
0.0713,
0.0048,
0.0402,
0.0071,
0.0251,
-0.0227,
-0.0367,
0.0651,
-0.1552,
0.0851,
-0.1552,
-0.1552,
-0.1552,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.0227,
-0.0367,
-0.0148,
-0.065,
0.0085,
-0.0337,
0.0713,
0.027,
-0.1454,
-0.0148,
0.0651,
-0.1552,
0.0851,
-0.1552,
-0.1552,
-0.1552,
-0.0058,
-0.0132,
-0.0004,
-0.001,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.1035,
0.3185,
-0.1353,
-0.1353,
0.0048,
0.0402,
-0.0227,
-0.0367,
-0.0148,
0.027,
-0.1454,
0.0285,
-0.1535,
0.0071,
0.0251,
0.0071,
0.0251,
0.0071,
0.0251,
-0.0148,
0.0307,
-0.0772,
-0.0227,
-0.0367,
-0.1035,
0.3185,
-0.1353,
-0.1353,
0.0044,
0.0249,
0.0071,
0.0251,
0.0085,
-0.0337,
0.0713,
0.027,
-0.1454,
-0.0148,
-0.065,
-0.0148,
-0.065,
0.0369,
-0.1135,
-0.088,
-0.088,
-0.0148,
-0.0148,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.0004,
-0.001,
0.0231,
-0.1155,
0.0071,
0.0251,
0.0307,
-0.0772,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
0.0231,
-0.1155,
-0.0148,
0.0369,
-0.1135,
-0.088,
-0.088,
0.0044,
0.0249,
0.0209,
-0.1029,
-0.0148,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
0.0048,
0.0402,
0.0651,
-0.1552,
0.0851,
-0.1552,
-0.1552,
-0.1552,
0.027,
-0.1454,
-0.0148,
0.0052,
0.0006,
0.0436,
0.0209,
-0.1029,
0.0307,
-0.0772,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
0.0085,
-0.0337,
0.0713,
-0.0148,
-0.0058,
-0.0132,
0.0231,
-0.1155,
0.0044,
0.0249,
0.0071,
0.0251,
-0.0148,
-0.065,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
0.0085,
-0.0337,
0.0713,
-0.065,
-0.0004,
-0.001,
-0.0148,
0.0231,
-0.1155,
-0.0004,
-0.001,
0.027,
-0.1454,
-0.0227,
-0.0367,
-0.065,
0.0085,
-0.0337,
0.0713,
0.027,
-0.1454,
-0.0148,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
0.0307,
-0.0772,
0.0285,
-0.1535,
-0.0227,
-0.0367,
0.0048,
0.0402,
0.0048,
0.0402,
0.027,
-0.1454,
0.0048,
0.0402,
0.0285,
-0.1535,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.0227,
-0.0367,
0.0052,
0.0006,
0.0436,
0.027,
-0.1454,
-0.0148,
-0.0148,
0.0209,
-0.1029,
0.0231,
-0.1155,
0.0651,
-0.1552,
0.0851,
-0.1552,
-0.1552,
-0.1552,
0.0052,
0.0006,
0.0436,
-0.065,
0.0048,
0.0402,
-0.0227,
-0.0367,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.0058,
-0.0132,
0.0071,
0.0251,
0.0231,
-0.1155,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.0148,
0.0085,
-0.0337,
0.0713,
0.0071,
0.0251,
-0.1035,
0.3185,
-0.1353,
-0.1353,
0.0048,
0.0402,
-0.0227,
-0.0367,
-0.0148,
0.0231,
-0.1155,
-0.0058,
-0.0132,
0.0307,
-0.0772,
0.0231,
-0.1155,
0.0369,
-0.1135,
-0.088,
-0.088,
-0.065,
-0.0148,
-0.0148,
0.0231,
-0.1155,
0.0044,
0.0249,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.065,
0.0285,
-0.1535,
-0.0227,
-0.0367,
0.0307,
-0.0772,
0.0044,
0.0249,
0.0285,
-0.1535,
-0.065,
-0.0227,
-0.0367,
0.0052,
0.0006,
0.0436,
0.027,
-0.1454,
0.0044,
0.0249,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
-0.0004,
-0.001,
0.0651,
-0.1552,
0.0851,
-0.1552,
-0.1552,
-0.1552,
-0.0227,
-0.0367,
0.0071,
0.0251,
0.0071,
0.0251,
0.0285,
-0.1535,
-0.0148,
0.0048,
0.0402,
-0.065,
-0.1035,
0.3185,
-0.1353,
-0.1353,
-0.0227,
-0.0367,
0.0285,
-0.1535,
-0.0148,
-0.0227,
-0.0367,
0.0052,
0.0006,
0.0436,
0.0307,
-0.0772,
0.0048,
0.0402,
0.0071,
0.0251,
-0.0148,
0.0209,
-0.1029,
0.027,
-0.1454,
-0.0058,
-0.0132,
0.027,
-0.1454,
-0.0148,
0.0231,
-0.1155,
-0.0058,
-0.0132,
0.0607,
-0.1868,
-0.1447,
-0.1447,
0.1377,
0.0052,
0.0006,
0.0436,
0.0369,
-0.1135,
-0.088,
-0.088,
-0.0148;
	particlenames = 
"MBB",
"MSC1",
"ABB",
"PBB",
"PSC1",
"KBB",
"KSC1",
"KSC2",
"DBB",
"DSC1",
"NBB",
"NSC1",
"TBB",
"TSC1",
"WBB",
"WSC1",
"WSC2",
"WSC3",
"WSC4",
"WSC5",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"TBB",
"TSC1",
"GBB",
"ABB",
"KBB",
"KSC1",
"KSC2",
"LBB",
"LSC1",
"GBB",
"WBB",
"WSC1",
"WSC2",
"WSC3",
"WSC4",
"WSC5",
"SBB",
"SSC1",
"QBB",
"QSC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"HBB",
"HSC1",
"HSC2",
"HSC3",
"DBB",
"DSC1",
"TBB",
"TSC1",
"GBB",
"LBB",
"LSC1",
"IBB",
"ISC1",
"NBB",
"NSC1",
"NBB",
"NSC1",
"NBB",
"NSC1",
"GBB",
"PBB",
"PSC1",
"TBB",
"TSC1",
"HBB",
"HSC1",
"HSC2",
"HSC3",
"EBB",
"ESC1",
"NBB",
"NSC1",
"KBB",
"KSC1",
"KSC2",
"LBB",
"LSC1",
"GBB",
"ABB",
"GBB",
"ABB",
"FBB",
"FSC1",
"FSC2",
"FSC3",
"GBB",
"GBB",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"QBB",
"QSC1",
"VBB",
"VSC1",
"NBB",
"NSC1",
"PBB",
"PSC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"VBB",
"VSC1",
"GBB",
"FBB",
"FSC1",
"FSC2",
"FSC3",
"EBB",
"ESC1",
"MBB",
"MSC1",
"GBB",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"DBB",
"DSC1",
"WBB",
"WSC1",
"WSC2",
"WSC3",
"WSC4",
"WSC5",
"LBB",
"LSC1",
"GBB",
"RBB",
"RSC1",
"RSC2",
"MBB",
"MSC1",
"PBB",
"PSC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"KBB",
"KSC1",
"KSC2",
"GBB",
"SBB",
"SSC1",
"VBB",
"VSC1",
"EBB",
"ESC1",
"NBB",
"NSC1",
"GBB",
"ABB",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"KBB",
"KSC1",
"KSC2",
"ABB",
"QBB",
"QSC1",
"GBB",
"VBB",
"VSC1",
"QBB",
"QSC1",
"LBB",
"LSC1",
"TBB",
"TSC1",
"ABB",
"KBB",
"KSC1",
"KSC2",
"LBB",
"LSC1",
"GBB",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"PBB",
"PSC1",
"IBB",
"ISC1",
"TBB",
"TSC1",
"DBB",
"DSC1",
"DBB",
"DSC1",
"LBB",
"LSC1",
"DBB",
"DSC1",
"IBB",
"ISC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"TBB",
"TSC1",
"RBB",
"RSC1",
"RSC2",
"LBB",
"LSC1",
"GBB",
"GBB",
"MBB",
"MSC1",
"VBB",
"VSC1",
"WBB",
"WSC1",
"WSC2",
"WSC3",
"WSC4",
"WSC5",
"RBB",
"RSC1",
"RSC2",
"ABB",
"DBB",
"DSC1",
"TBB",
"TSC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"SBB",
"SSC1",
"NBB",
"NSC1",
"VBB",
"VSC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"GBB",
"KBB",
"KSC1",
"KSC2",
"NBB",
"NSC1",
"HBB",
"HSC1",
"HSC2",
"HSC3",
"DBB",
"DSC1",
"TBB",
"TSC1",
"GBB",
"VBB",
"VSC1",
"SBB",
"SSC1",
"PBB",
"PSC1",
"VBB",
"VSC1",
"FBB",
"FSC1",
"FSC2",
"FSC3",
"ABB",
"GBB",
"GBB",
"VBB",
"VSC1",
"EBB",
"ESC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"ABB",
"IBB",
"ISC1",
"TBB",
"TSC1",
"PBB",
"PSC1",
"EBB",
"ESC1",
"IBB",
"ISC1",
"ABB",
"TBB",
"TSC1",
"RBB",
"RSC1",
"RSC2",
"LBB",
"LSC1",
"EBB",
"ESC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"QBB",
"QSC1",
"WBB",
"WSC1",
"WSC2",
"WSC3",
"WSC4",
"WSC5",
"TBB",
"TSC1",
"NBB",
"NSC1",
"NBB",
"NSC1",
"IBB",
"ISC1",
"GBB",
"DBB",
"DSC1",
"ABB",
"HBB",
"HSC1",
"HSC2",
"HSC3",
"TBB",
"TSC1",
"IBB",
"ISC1",
"GBB",
"TBB",
"TSC1",
"RBB",
"RSC1",
"RSC2",
"PBB",
"PSC1",
"DBB",
"DSC1",
"NBB",
"NSC1",
"GBB",
"MBB",
"MSC1",
"LBB",
"LSC1",
"SBB",
"SSC1",
"LBB",
"LSC1",
"GBB",
"VBB",
"VSC1",
"SBB",
"SSC1",
"YBB",
"YSC1",
"YSC2",
"YSC3",
"YSC4",
"RBB",
"RSC1",
"RSC2",
"FBB",
"FSC1",
"FSC2",
"FSC3",
"GBB";
	resnames = 
"MET",
"MET",
"ALA",
"PRO",
"PRO",
"LYS",
"LYS",
"LYS",
"ASP",
"ASP",
"ASN",
"ASN",
"THR",
"THR",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"THR",
"THR",
"GLY",
"ALA",
"LYS",
"LYS",
"LYS",
"LEU",
"LEU",
"GLY",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"SER",
"SER",
"GLN",
"GLN",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"HIS",
"HIS",
"HIS",
"HIS",
"ASP",
"ASP",
"THR",
"THR",
"GLY",
"LEU",
"LEU",
"ILE",
"ILE",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"GLY",
"PRO",
"PRO",
"THR",
"THR",
"HIS",
"HIS",
"HIS",
"HIS",
"GLU",
"GLU",
"ASN",
"ASN",
"LYS",
"LYS",
"LYS",
"LEU",
"LEU",
"GLY",
"ALA",
"GLY",
"ALA",
"PHE",
"PHE",
"PHE",
"PHE",
"GLY",
"GLY",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"GLN",
"GLN",
"VAL",
"VAL",
"ASN",
"ASN",
"PRO",
"PRO",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"VAL",
"VAL",
"GLY",
"PHE",
"PHE",
"PHE",
"PHE",
"GLU",
"GLU",
"MET",
"MET",
"GLY",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"ASP",
"ASP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"LEU",
"LEU",
"GLY",
"ARG",
"ARG",
"ARG",
"MET",
"MET",
"PRO",
"PRO",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"LYS",
"LYS",
"LYS",
"GLY",
"SER",
"SER",
"VAL",
"VAL",
"GLU",
"GLU",
"ASN",
"ASN",
"GLY",
"ALA",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"LYS",
"LYS",
"LYS",
"ALA",
"GLN",
"GLN",
"GLY",
"VAL",
"VAL",
"GLN",
"GLN",
"LEU",
"LEU",
"THR",
"THR",
"ALA",
"LYS",
"LYS",
"LYS",
"LEU",
"LEU",
"GLY",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"PRO",
"PRO",
"ILE",
"ILE",
"THR",
"THR",
"ASP",
"ASP",
"ASP",
"ASP",
"LEU",
"LEU",
"ASP",
"ASP",
"ILE",
"ILE",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"THR",
"THR",
"ARG",
"ARG",
"ARG",
"LEU",
"LEU",
"GLY",
"GLY",
"MET",
"MET",
"VAL",
"VAL",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"ARG",
"ARG",
"ARG",
"ALA",
"ASP",
"ASP",
"THR",
"THR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"SER",
"SER",
"ASN",
"ASN",
"VAL",
"VAL",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"GLY",
"LYS",
"LYS",
"LYS",
"ASN",
"ASN",
"HIS",
"HIS",
"HIS",
"HIS",
"ASP",
"ASP",
"THR",
"THR",
"GLY",
"VAL",
"VAL",
"SER",
"SER",
"PRO",
"PRO",
"VAL",
"VAL",
"PHE",
"PHE",
"PHE",
"PHE",
"ALA",
"GLY",
"GLY",
"VAL",
"VAL",
"GLU",
"GLU",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"ALA",
"ILE",
"ILE",
"THR",
"THR",
"PRO",
"PRO",
"GLU",
"GLU",
"ILE",
"ILE",
"ALA",
"THR",
"THR",
"ARG",
"ARG",
"ARG",
"LEU",
"LEU",
"GLU",
"GLU",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"GLN",
"GLN",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"THR",
"THR",
"ASN",
"ASN",
"ASN",
"ASN",
"ILE",
"ILE",
"GLY",
"ASP",
"ASP",
"ALA",
"HIS",
"HIS",
"HIS",
"HIS",
"THR",
"THR",
"ILE",
"ILE",
"GLY",
"THR",
"THR",
"ARG",
"ARG",
"ARG",
"PRO",
"PRO",
"ASP",
"ASP",
"ASN",
"ASN",
"GLY",
"MET",
"MET",
"LEU",
"LEU",
"SER",
"SER",
"LEU",
"LEU",
"GLY",
"VAL",
"VAL",
"SER",
"SER",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"ARG",
"ARG",
"ARG",
"PHE",
"PHE",
"PHE",
"PHE",
"GLY";
	resids = 
0,
0,
1,
2,
2,
3,
3,
3,
4,
4,
5,
5,
6,
6,
7,
7,
7,
7,
7,
7,
8,
8,
8,
8,
8,
9,
9,
10,
11,
12,
12,
12,
13,
13,
14,
15,
15,
15,
15,
15,
15,
16,
16,
17,
17,
18,
18,
18,
18,
18,
19,
19,
19,
19,
20,
20,
21,
21,
22,
23,
23,
24,
24,
25,
25,
26,
26,
27,
27,
28,
29,
29,
30,
30,
31,
31,
31,
31,
32,
32,
33,
33,
34,
34,
34,
35,
35,
36,
37,
38,
39,
40,
40,
40,
40,
41,
42,
43,
43,
43,
43,
43,
44,
44,
45,
45,
46,
46,
47,
47,
48,
48,
48,
48,
48,
49,
49,
50,
51,
51,
51,
51,
52,
52,
53,
53,
54,
55,
55,
55,
55,
55,
56,
56,
57,
57,
57,
57,
57,
57,
58,
58,
59,
60,
60,
60,
61,
61,
62,
62,
63,
63,
63,
63,
63,
64,
64,
64,
65,
66,
66,
67,
67,
68,
68,
69,
69,
70,
71,
72,
72,
72,
72,
72,
73,
73,
73,
74,
75,
75,
76,
77,
77,
78,
78,
79,
79,
80,
80,
81,
82,
82,
82,
83,
83,
84,
85,
85,
85,
85,
85,
86,
86,
87,
87,
88,
88,
89,
89,
90,
90,
91,
91,
92,
92,
93,
93,
94,
94,
94,
94,
94,
95,
95,
96,
96,
96,
97,
97,
98,
99,
100,
100,
101,
101,
102,
102,
102,
102,
102,
102,
103,
103,
103,
104,
105,
105,
106,
106,
107,
107,
107,
107,
107,
108,
108,
109,
109,
110,
110,
111,
111,
111,
111,
111,
112,
113,
113,
113,
114,
114,
115,
115,
115,
115,
116,
116,
117,
117,
118,
119,
119,
120,
120,
121,
121,
122,
122,
123,
123,
123,
123,
124,
125,
126,
127,
127,
128,
128,
129,
129,
129,
129,
129,
130,
131,
131,
132,
132,
133,
133,
134,
134,
135,
135,
136,
137,
137,
138,
138,
138,
139,
139,
140,
140,
141,
141,
141,
141,
141,
142,
142,
143,
143,
143,
143,
143,
143,
144,
144,
145,
145,
146,
146,
147,
147,
148,
149,
149,
150,
151,
151,
151,
151,
152,
152,
153,
153,
154,
155,
155,
156,
156,
156,
157,
157,
158,
158,
159,
159,
160,
161,
161,
162,
162,
163,
163,
164,
164,
165,
166,
166,
167,
167,
168,
168,
168,
168,
168,
169,
169,
169,
170,
170,
170,
170,
171;
	chainnames = 
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A";
	dynamicstate = 
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1;
	nbspringsperparticle = 
5,
1,
4,
5,
6,
4,
2,
1,
7,
2,
6,
3,
8,
6,
10,
7,
7,
7,
6,
6,
9,
9,
9,
9,
7,
8,
4,
7,
5,
6,
7,
4,
6,
2,
5,
8,
7,
6,
7,
7,
5,
6,
9,
7,
1,
9,
6,
5,
5,
4,
8,
8,
6,
7,
6,
6,
4,
2,
3,
3,
2,
4,
2,
4,
2,
6,
3,
3,
2,
3,
4,
3,
5,
4,
6,
4,
3,
4,
5,
4,
5,
2,
5,
8,
7,
5,
2,
3,
9,
5,
4,
6,
7,
7,
8,
4,
9,
8,
10,
10,
6,
5,
9,
6,
6,
3,
8,
8,
7,
4,
9,
7,
7,
6,
3,
7,
4,
8,
6,
4,
5,
4,
5,
6,
4,
1,
5,
7,
6,
7,
6,
7,
9,
3,
7,
10,
8,
6,
8,
5,
6,
4,
4,
4,
4,
3,
6,
2,
5,
3,
5,
5,
6,
5,
3,
4,
4,
2,
4,
4,
3,
5,
3,
4,
3,
3,
4,
3,
4,
6,
7,
6,
7,
4,
7,
2,
3,
3,
4,
3,
6,
5,
3,
5,
5,
5,
2,
6,
7,
5,
5,
8,
2,
6,
2,
5,
8,
7,
7,
6,
3,
8,
6,
5,
3,
6,
5,
5,
1,
7,
4,
7,
5,
6,
4,
5,
2,
7,
9,
8,
7,
8,
7,
3,
6,
7,
5,
6,
2,
4,
4,
5,
6,
6,
2,
7,
8,
8,
7,
11,
7,
6,
4,
4,
6,
5,
5,
5,
5,
8,
7,
7,
5,
4,
10,
8,
5,
2,
5,
6,
7,
8,
5,
6,
4,
6,
3,
3,
1,
6,
2,
6,
7,
4,
4,
8,
4,
7,
3,
10,
5,
2,
5,
7,
5,
3,
7,
7,
8,
7,
3,
5,
6,
3,
8,
6,
5,
6,
4,
8,
7,
7,
5,
4,
7,
5,
2,
7,
6,
6,
4,
9,
3,
6,
3,
7,
5,
4,
5,
6,
6,
4,
2,
7,
4,
8,
7,
8,
8,
5,
9,
4,
8,
9,
8,
8,
10,
6,
6,
6,
5,
2,
4,
5,
6,
1,
4,
3,
2,
5,
6,
7,
6,
9,
7,
6,
7,
2,
5,
5,
3,
4,
7,
5,
3,
4,
4,
6,
8,
5,
7,
5,
3,
8,
5,
5,
7,
5,
2,
5,
5,
3,
6,
8,
8,
6,
6,
8,
4,
9,
6,
5,
5,
6,
3,
6,
2;
	springs = 
0, 1,
0, 2,
2, 3,
3, 4,
3, 5,
5, 6,
5, 8,
6, 7,
8, 9,
8, 10,
10, 11,
10, 12,
12, 13,
12, 14,
14, 15,
14, 20,
15, 16,
15, 18,
16, 19,
18, 19,
20, 21,
20, 25,
21, 22,
21, 23,
22, 23,
22, 24,
23, 24,
25, 26,
25, 27,
27, 28,
28, 29,
29, 30,
29, 32,
30, 31,
32, 33,
32, 34,
34, 35,
35, 36,
35, 41,
36, 37,
36, 39,
37, 40,
39, 40,
41, 42,
41, 43,
43, 44,
43, 45,
45, 46,
45, 50,
46, 47,
46, 48,
47, 48,
47, 49,
48, 49,
50, 51,
50, 54,
51, 52,
51, 53,
52, 53,
54, 55,
54, 56,
56, 57,
56, 58,
58, 59,
59, 60,
59, 61,
61, 62,
61, 63,
61, 65,
63, 64,
63, 65,
65, 66,
65, 67,
67, 68,
67, 69,
69, 70,
70, 71,
70, 72,
72, 73,
72, 74,
74, 75,
74, 78,
75, 76,
75, 77,
76, 77,
78, 79,
78, 80,
80, 81,
80, 82,
82, 83,
82, 85,
83, 84,
85, 86,
85, 87,
87, 88,
88, 89,
89, 90,
90, 91,
91, 92,
91, 95,
92, 93,
92, 94,
93, 94,
95, 96,
96, 97,
97, 98,
97, 102,
98, 99,
98, 100,
99, 100,
99, 101,
100, 101,
102, 103,
102, 104,
104, 105,
104, 106,
106, 107,
106, 108,
108, 109,
108, 110,
110, 111,
110, 115,
111, 112,
111, 113,
112, 113,
112, 114,
113, 114,
115, 116,
115, 117,
117, 118,
118, 119,
118, 122,
119, 120,
119, 121,
120, 121,
122, 123,
122, 124,
124, 125,
124, 126,
126, 127,
127, 128,
127, 132,
128, 129,
128, 130,
129, 130,
129, 131,
130, 131,
132, 133,
132, 134,
134, 135,
134, 140,
135, 136,
135, 138,
136, 139,
138, 139,
140, 141,
140, 142,
142, 143,
143, 144,
143, 146,
144, 145,
146, 147,
146, 148,
148, 149,
148, 150,
150, 151,
150, 155,
151, 152,
151, 153,
152, 153,
152, 154,
153, 154,
155, 156,
156, 157,
158, 159,
159, 160,
159, 161,
161, 162,
161, 163,
161, 164,
162, 164,
163, 164,
165, 166,
165, 167,
167, 168,
168, 169,
169, 170,
169, 174,
170, 171,
170, 172,
171, 172,
171, 173,
172, 173,
174, 175,
174, 177,
175, 176,
177, 178,
178, 179,
178, 180,
180, 181,
181, 182,
181, 183,
183, 184,
183, 185,
185, 186,
185, 187,
187, 188,
187, 189,
189, 190,
190, 191,
190, 193,
191, 192,
193, 194,
193, 195,
195, 196,
196, 197,
196, 201,
197, 198,
197, 199,
198, 199,
198, 200,
199, 200,
201, 202,
201, 203,
203, 204,
203, 205,
205, 206,
205, 207,
207, 208,
207, 209,
209, 210,
209, 211,
211, 212,
211, 213,
213, 214,
213, 215,
215, 216,
215, 217,
217, 218,
217, 222,
218, 219,
218, 220,
219, 220,
219, 221,
220, 221,
222, 223,
222, 224,
224, 225,
224, 227,
225, 226,
227, 228,
227, 229,
229, 230,
230, 231,
231, 232,
231, 233,
233, 234,
233, 235,
235, 236,
235, 241,
236, 237,
236, 239,
237, 240,
239, 240,
241, 242,
241, 244,
242, 243,
244, 245,
245, 246,
245, 247,
247, 248,
247, 249,
249, 250,
249, 254,
250, 251,
250, 252,
251, 252,
251, 253,
252, 253,
254, 255,
254, 256,
256, 257,
256, 258,
258, 259,
258, 260,
260, 261,
260, 265,
261, 262,
261, 263,
262, 263,
262, 264,
263, 264,
265, 266,
266, 267,
266, 269,
267, 268,
269, 270,
269, 271,
271, 272,
271, 275,
272, 273,
272, 274,
273, 274,
275, 276,
275, 277,
277, 278,
277, 279,
279, 280,
280, 281,
280, 282,
282, 283,
282, 284,
284, 285,
284, 286,
286, 287,
286, 288,
288, 289,
288, 292,
289, 290,
289, 291,
290, 291,
292, 293,
293, 294,
294, 295,
295, 296,
295, 297,
297, 298,
297, 299,
299, 300,
299, 304,
300, 301,
300, 302,
301, 302,
301, 303,
302, 303,
304, 305,
305, 306,
305, 307,
307, 308,
307, 309,
309, 310,
309, 311,
311, 312,
311, 313,
313, 314,
313, 315,
315, 316,
316, 317,
316, 318,
318, 319,
318, 321,
319, 320,
321, 322,
321, 323,
323, 324,
323, 325,
325, 326,
325, 330,
326, 327,
326, 328,
327, 328,
327, 329,
328, 329,
330, 331,
330, 332,
332, 333,
332, 338,
333, 334,
333, 336,
334, 337,
336, 337,
338, 339,
338, 340,
340, 341,
340, 342,
342, 343,
344, 345,
344, 346,
346, 347,
347, 348,
347, 349,
349, 350,
350, 351,
350, 354,
351, 352,
351, 353,
351, 354,
351, 355,
352, 353,
352, 355,
353, 354,
354, 355,
354, 356,
356, 357,
356, 358,
358, 359,
358, 363,
359, 360,
359, 361,
359, 362,
361, 362,
361, 364,
361, 365,
362, 363,
364, 365,
364, 366,
366, 367,
366, 368,
368, 369,
368, 370,
370, 371,
371, 372,
371, 373,
373, 374,
373, 375,
375, 376,
375, 377,
377, 378,
377, 379,
379, 380,
380, 381,
380, 382,
382, 383,
382, 384,
384, 385,
384, 389,
385, 386,
385, 387,
386, 387,
386, 388,
387, 388,
389, 390,
389, 392,
390, 391,
392, 393,
392, 396,
393, 394,
393, 395,
394, 395,
0, 209,
0, 214,
0, 391,
2, 4,
2, 391,
3, 391,
3, 103,
4, 390,
4, 391,
4, 103,
4, 22,
5, 13,
8, 13,
8, 104,
8, 11,
8, 102,
9, 106,
10, 13,
10, 99,
10, 101,
11, 101,
12, 15,
12, 102,
12, 98,
12, 16,
12, 99,
13, 396,
13, 14,
14, 21,
14, 22,
14, 392,
14, 393,
14, 16,
14, 17,
15, 20,
15, 17,
15, 19,
16, 99,
16, 17,
16, 18,
17, 98,
17, 99,
17, 18,
17, 19,
18, 96,
18, 98,
19, 98,
19, 99,
20, 26,
20, 395,
20, 22,
20, 23,
20, 96,
21, 390,
21, 383,
21, 25,
21, 24,
21, 96,
22, 103,
22, 96,
22, 97,
23, 383,
23, 94,
23, 25,
23, 123,
23, 96,
24, 192,
24, 123,
24, 96,
24, 97,
25, 383,
25, 94,
25, 384,
26, 27,
26, 395,
27, 93,
27, 94,
27, 91,
27, 92,
28, 30,
28, 380,
28, 93,
29, 33,
29, 89,
29, 88,
30, 32,
30, 376,
30, 89,
30, 93,
31, 376,
31, 331,
31, 133,
32, 377,
32, 376,
34, 36,
34, 39,
34, 87,
35, 37,
35, 38,
35, 39,
35, 373,
35, 42,
36, 38,
36, 40,
36, 41,
37, 38,
37, 374,
37, 39,
38, 40,
38, 374,
38, 39,
38, 373,
39, 373,
40, 374,
41, 82,
41, 83,
42, 43,
42, 53,
42, 370,
42, 45,
42, 51,
42, 83,
42, 52,
43, 48,
43, 78,
43, 46,
45, 48,
45, 47,
45, 369,
45, 51,
45, 54,
46, 49,
46, 54,
47, 369,
49, 369,
50, 53,
50, 84,
50, 55,
50, 52,
50, 368,
51, 83,
51, 84,
51, 368,
52, 368,
52, 367,
53, 370,
53, 368,
53, 367,
54, 57,
55, 79,
55, 56,
55, 84,
55, 172,
58, 60,
62, 65,
63, 66,
64, 66,
65, 68,
69, 71,
70, 73,
71, 166,
72, 77,
72, 75,
73, 74,
73, 155,
74, 76,
74, 77,
78, 81,
79, 84,
79, 145,
80, 146,
80, 83,
82, 86,
83, 141,
83, 142,
84, 171,
84, 173,
85, 141,
85, 142,
88, 134,
88, 137,
88, 138,
88, 139,
88, 135,
88, 136,
89, 138,
90, 92,
90, 127,
91, 93,
91, 94,
92, 123,
92, 95,
93, 320,
94, 383,
94, 320,
95, 124,
96, 98,
97, 100,
97, 118,
97, 99,
98, 102,
98, 101,
99, 102,
100, 102,
100, 105,
102, 105,
103, 106,
103, 115,
104, 107,
104, 115,
106, 109,
106, 110,
106, 115,
107, 109,
107, 108,
107, 110,
107, 111,
107, 116,
107, 115,
108, 112,
108, 111,
108, 113,
109, 113,
110, 112,
110, 195,
110, 113,
110, 116,
111, 114,
111, 195,
112, 202,
112, 198,
116, 117,
117, 190,
117, 191,
117, 119,
117, 121,
117, 120,
118, 121,
118, 120,
120, 189,
122, 188,
122, 187,
123, 320,
123, 191,
126, 184,
126, 128,
126, 183,
127, 133,
127, 130,
127, 129,
128, 132,
128, 131,
129, 132,
129, 179,
129, 180,
130, 138,
130, 132,
131, 138,
131, 135,
131, 132,
131, 179,
132, 135,
132, 180,
134, 141,
134, 137,
134, 136,
135, 140,
135, 137,
135, 139,
135, 176,
136, 140,
136, 137,
136, 138,
136, 176,
137, 138,
137, 139,
140, 177,
143, 169,
144, 146,
144, 170,
145, 170,
146, 149,
147, 149,
148, 151,
148, 153,
150, 152,
150, 153,
151, 154,
152, 156,
152, 157,
155, 158,
156, 158,
158, 160,
159, 162,
160, 161,
163, 166,
163, 165,
166, 167,
168, 249,
168, 250,
169, 171,
169, 172,
170, 173,
170, 174,
171, 174,
172, 174,
172, 248,
174, 245,
178, 241,
180, 232,
180, 182,
181, 232,
181, 233,
182, 183,
184, 226,
184, 287,
184, 232,
185, 188,
185, 230,
186, 187,
187, 227,
188, 225,
188, 226,
188, 189,
188, 227,
189, 227,
190, 194,
191, 218,
191, 219,
191, 193,
191, 225,
193, 218,
193, 222,
195, 197,
196, 199,
196, 202,
196, 214,
196, 215,
196, 198,
197, 200,
197, 201,
197, 202,
198, 201,
198, 202,
199, 201,
199, 202,
201, 204,
201, 205,
203, 206,
203, 211,
204, 216,
205, 209,
205, 211,
206, 207,
206, 209,
206, 211,
207, 210,
209, 304,
210, 303,
210, 304,
211, 214,
212, 302,
212, 300,
212, 213,
212, 296,
213, 296,
213, 297,
215, 218,
217, 294,
217, 219,
217, 220,
217, 223,
218, 294,
218, 221,
218, 222,
219, 294,
219, 222,
219, 225,
220, 294,
220, 295,
220, 298,
221, 294,
221, 295,
221, 319,
221, 324,
221, 320,
222, 225,
223, 224,
224, 292,
224, 228,
225, 292,
226, 324,
226, 331,
229, 286,
229, 287,
230, 287,
231, 282,
231, 234,
232, 287,
232, 233,
233, 236,
235, 237,
235, 238,
235, 239,
235, 279,
236, 238,
236, 240,
236, 241,
236, 279,
237, 238,
237, 239,
237, 283,
237, 279,
237, 280,
238, 239,
238, 240,
238, 279,
238, 277,
239, 276,
239, 241,
239, 244,
239, 275,
239, 279,
239, 277,
240, 276,
240, 279,
240, 277,
242, 246,
242, 244,
243, 246,
243, 272,
243, 274,
244, 246,
244, 275,
245, 248,
246, 272,
247, 250,
247, 269,
248, 249,
248, 269,
249, 255,
249, 251,
249, 252,
250, 254,
250, 253,
251, 254,
251, 265,
251, 267,
252, 254,
253, 254,
254, 257,
254, 260,
254, 265,
255, 256,
255, 258,
255, 261,
255, 263,
255, 260,
255, 265,
256, 259,
258, 261,
259, 261,
259, 262,
259, 263,
259, 264,
260, 262,
260, 263,
261, 264,
261, 265,
269, 272,
270, 271,
271, 273,
271, 274,
272, 275,
273, 275,
275, 278,
276, 277,
278, 279,
279, 281,
280, 283,
282, 285,
283, 339,
283, 343,
283, 285,
283, 284,
284, 287,
286, 289,
286, 291,
286, 290,
287, 288,
288, 332,
288, 335,
288, 336,
288, 337,
289, 335,
289, 337,
289, 334,
291, 334,
291, 341,
292, 325,
292, 336,
293, 325,
294, 296,
295, 321,
296, 297,
297, 300,
298, 319,
298, 320,
299, 301,
299, 302,
299, 317,
299, 315,
299, 316,
300, 303,
300, 304,
301, 305,
301, 306,
301, 304,
304, 307,
305, 308,
307, 310,
307, 313,
307, 311,
308, 309,
308, 310,
308, 313,
308, 311,
309, 313,
309, 312,
310, 312,
311, 314,
311, 386,
311, 390,
311, 389,
314, 315,
315, 317,
315, 382,
315, 383,
316, 319,
317, 318,
318, 379,
319, 379,
322, 323,
323, 326,
323, 375,
323, 376,
324, 325,
325, 327,
325, 328,
326, 329,
326, 336,
326, 330,
327, 374,
327, 371,
327, 370,
327, 330,
328, 335,
328, 336,
328, 333,
328, 330,
329, 370,
329, 333,
330, 371,
330, 336,
330, 333,
331, 372,
332, 335,
332, 336,
332, 334,
332, 339,
333, 335,
333, 337,
333, 338,
334, 335,
334, 336,
334, 338,
335, 336,
335, 337,
338, 367,
339, 367,
339, 340,
339, 343,
340, 343,
342, 362,
342, 344,
343, 344,
344, 362,
344, 363,
346, 363,
346, 348,
349, 353,
349, 351,
349, 354,
350, 353,
350, 352,
350, 355,
351, 356,
352, 356,
352, 354,
353, 356,
353, 357,
353, 358,
353, 355,
355, 356,
358, 360,
359, 363,
360, 362,
362, 365,
365, 366,
367, 368,
369, 370,
372, 373,
373, 376,
375, 378,
376, 377,
379, 381,
380, 383,
381, 382,
382, 385,
383, 384,
384, 386,
384, 390,
384, 387,
385, 388,
385, 389,
386, 389,
387, 389,
387, 394,
387, 395,
387, 393,
388, 389,
389, 393,
392, 395;
	springsstiffness = 
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30;
	springsequilibrium = 
3.49113,
3.2253,
3.04695,
2.39325,
3.22338,
3.38844,
3.31428,
2.89512,
3.12214,
3.57116,
3.13078,
3.36313,
2.59595,
3.48745,
2.66662,
3.66438,
2.40212,
3.4954,
3.52986,
2.12387,
2.40836,
3.6637,
2.46271,
2.49497,
2.40557,
2.3754,
2.397,
2.55297,
3.72952,
3.59985,
3.72721,
3.03653,
3.53875,
3.18502,
3.37071,
3.5208,
3.68383,
2.39598,
3.60453,
2.40717,
3.52645,
3.52576,
2.12533,
2.44589,
3.60134,
2.97177,
3.22161,
2.36338,
3.65997,
2.46797,
2.47586,
2.38803,
2.38484,
2.38352,
2.52165,
3.1871,
2.38786,
2.36632,
1.74536,
2.9429,
3.74665,
2.75813,
3.72715,
3.62383,
3.42398,
3.87543,
3.18712,
2.26768,
3.06026,
3.44322,
2.86216,
3.2124,
3.22599,
3.2838,
3.71923,
3.17701,
2.2621,
3.73344,
2.50777,
3.23825,
2.87498,
3.80048,
2.07075,
2.07033,
1.79016,
3.83325,
3.7016,
3.27337,
3.59278,
3.08951,
3.55738,
2.69522,
3.37186,
3.70837,
3.54218,
3.7159,
3.62933,
3.70993,
2.54612,
3.61143,
2.39963,
2.41088,
1.85542,
3.71817,
3.6196,
2.52858,
3.3929,
2.46843,
2.46817,
2.39394,
2.38932,
2.3811,
3.62372,
3.53979,
2.59008,
3.15455,
2.78328,
3.47102,
2.4421,
3.3893,
2.57274,
3.38971,
2.45253,
2.47179,
2.40135,
2.38456,
2.40645,
2.51612,
3.60962,
3.60417,
2.9236,
3.69302,
2.38181,
2.37209,
1.84482,
3.91033,
3.52267,
3.77109,
3.65247,
3.58168,
2.48026,
3.58859,
2.4641,
2.46829,
2.40377,
2.38761,
2.37346,
3.3421,
3.66434,
2.4111,
3.65201,
2.3776,
3.54558,
3.54089,
2.10431,
3.45606,
3.59185,
3.20798,
3.02019,
3.48508,
2.98278,
3.53282,
3.40954,
2.16323,
3.80027,
2.50079,
3.19084,
2.47594,
2.4501,
2.38936,
2.38965,
2.3814,
3.41245,
3.1105,
3.62399,
2.04596,
2.82127,
2.43054,
3.52721,
2.90801,
2.91688,
3.81439,
3.28981,
3.44965,
3.56143,
3.81864,
2.48574,
3.60687,
2.48499,
2.48009,
2.39577,
2.39312,
2.40038,
3.16834,
3.59305,
2.85247,
3.64004,
3.95215,
3.77932,
3.53013,
2.51778,
3.59099,
3.74535,
3.69952,
3.08586,
3.62584,
2.59513,
3.47038,
3.66355,
3.09691,
3.58822,
2.75914,
3.34455,
3.62825,
3.64962,
2.50873,
3.46736,
2.46644,
2.45783,
2.40934,
2.38859,
2.38705,
2.0724,
3.43794,
2.66005,
3.13641,
2.65439,
3.55278,
3.204,
3.37791,
3.22098,
3.33818,
3.13773,
3.51425,
3.37299,
3.4707,
2.95784,
3.6521,
2.40524,
3.54141,
2.47547,
2.48533,
2.41829,
2.3932,
2.40777,
2.59354,
3.53877,
3.37092,
3.65301,
2.94105,
2.99587,
3.72747,
3.57753,
3.77238,
3.72558,
3.48396,
2.59945,
3.59456,
2.30993,
3.75096,
2.40269,
3.51025,
3.51214,
2.1354,
2.98399,
3.56411,
3.48958,
3.68762,
3.27695,
3.40737,
2.70311,
3.70667,
2.62003,
3.60626,
2.46684,
2.48171,
2.38979,
2.38267,
2.40125,
2.60676,
3.46889,
3.09249,
2.93706,
2.71444,
3.43434,
2.54755,
3.04266,
2.47317,
2.47726,
2.39511,
2.37269,
2.39124,
3.32583,
3.28562,
3.66521,
2.75413,
3.22993,
3.59406,
2.42483,
3.6419,
2.38814,
2.35119,
1.76424,
3.25104,
3.61262,
2.73831,
3.71658,
3.54636,
2.73144,
3.64464,
2.58188,
3.15314,
2.26383,
3.64494,
2.56371,
3.63435,
2.99637,
3.66099,
2.39535,
2.39819,
1.83075,
3.59967,
3.67166,
3.57121,
2.67537,
3.62012,
3.92663,
3.65379,
2.51179,
3.58732,
2.45624,
2.48208,
2.37731,
2.37918,
2.40772,
3.45297,
2.87104,
3.02379,
2.53641,
3.41271,
2.48692,
3.41483,
3.41999,
3.29864,
2.70881,
3.5785,
3.50073,
2.54146,
3.68736,
3.14085,
3.55872,
3.59784,
3.12195,
3.58025,
3.8542,
3.61192,
2.44974,
3.54048,
2.45686,
2.4847,
2.42503,
2.36366,
2.39655,
3.85335,
3.60432,
2.42886,
3.53131,
2.39958,
3.54636,
3.53688,
2.12685,
2.41312,
3.34095,
2.7459,
3.81789,
3.30384,
3.26788,
3.2231,
3.51905,
3.31969,
3.62411,
3.67084,
2.5001,
3.16445,
2.29529,
2.38633,
1.75726,
1.76447,
1.76771,
1.98854,
2.4226,
2.62861,
3.66902,
3.18273,
3.45918,
3.8885,
2.72702,
2.77663,
3.94922,
1.94869,
3.25735,
3.13562,
2.20926,
4.04597,
2.00075,
3.5892,
2.79183,
3.48357,
3.26435,
3.33731,
3.60812,
3.55499,
3.43274,
3.3489,
3.6992,
2.31854,
3.55376,
3.31878,
3.6139,
3.60756,
2.67268,
3.66528,
2.39455,
3.52435,
2.49544,
3.53436,
2.45833,
2.46388,
2.40999,
2.38124,
2.38981,
3.20564,
3.57267,
3.61445,
2.7966,
3.38694,
2.39952,
2.39716,
1.83818,
4.9487,
4.60654,
4.83631,
3.87331,
4.51582,
4.91516,
4.32741,
4.59717,
3.98261,
3.88723,
4.44996,
3.82807,
4.82775,
4.53438,
4.23386,
4.9593,
4.64987,
3.8805,
4.32467,
4.10135,
3.71242,
4.393,
4.27079,
4.99956,
4.57309,
3.94786,
4.28162,
4.47804,
4.27064,
4.80371,
4.57137,
4.83871,
4.56792,
4.87161,
4.75534,
2.43733,
4.46465,
4.02974,
1.81083,
3.86545,
4.25687,
4.06212,
2.07499,
2.07804,
4.25201,
4.16529,
4.20231,
4.40566,
4.35559,
4.55233,
4.04793,
3.96363,
3.98155,
4.94082,
4.94778,
4.43711,
4.2281,
4.6049,
4.99358,
3.75034,
4.33982,
4.85089,
4.44769,
4.98392,
4.83813,
4.26879,
4.16541,
3.86293,
4.14782,
4.76506,
4.31646,
4.97796,
3.98277,
4.75157,
4.3641,
3.71887,
4.04392,
3.84544,
4.3832,
4.956,
4.40503,
4.42818,
4.57563,
4.0375,
4.95071,
4.66319,
4.08166,
4.46967,
4.90222,
4.31619,
4.89163,
3.63676,
4.21251,
4.75165,
4.62703,
4.98108,
3.64534,
3.94221,
4.08972,
4.84725,
4.02032,
4.65468,
2.44759,
4.49251,
4.59623,
1.80218,
4.66085,
3.86181,
2.0923,
4.57922,
2.07702,
4.61032,
4.93316,
4.28114,
3.69577,
4.52141,
4.63047,
3.07743,
4.45992,
4.41693,
4.03765,
4.61206,
4.56656,
4.49643,
4.90113,
3.94045,
4.21391,
3.58628,
4.95943,
4.57112,
4.84169,
4.22803,
4.76991,
3.76111,
4.22915,
4.41274,
4.26387,
4.2017,
4.63412,
4.94258,
4.89271,
4.00309,
4.67649,
4.48758,
4.22948,
4.02208,
3.69368,
4.91388,
3.91034,
4.92405,
4.05411,
4.48911,
4.90004,
4.40386,
4.83245,
4.39687,
4.3137,
4.64873,
3.77033,
4.60485,
4.43981,
4.40994,
3.89696,
4.87963,
4.80137,
4.61371,
4.71699,
4.1842,
4.52746,
4.58347,
4.63496,
4.31814,
4.54371,
4.78445,
4.82982,
3.92326,
4.62055,
4.85837,
4.08151,
4.27133,
3.97444,
4.22243,
4.36414,
4.73464,
4.56842,
4.97934,
4.67134,
4.16732,
4.24879,
4.10523,
4.96487,
4.64614,
4.48721,
4.4566,
3.74037,
3.83883,
4.92509,
4.31018,
4.02843,
4.53876,
4.10062,
4.22177,
4.45761,
4.09739,
4.7942,
4.7873,
4.65342,
4.64974,
4.36644,
4.93862,
3.99221,
4.81526,
4.08189,
4.82149,
4.73375,
4.91081,
4.91474,
4.64403,
4.64695,
4.89016,
3.97942,
4.34432,
4.07251,
4.51028,
4.08523,
4.70882,
4.30388,
4.22227,
4.97358,
4.91807,
4.55529,
4.72716,
3.72628,
4.84513,
4.11198,
4.59359,
4.75013,
4.98281,
4.98711,
4.87488,
4.9882,
3.90383,
4.53376,
4.94073,
4.6685,
4.96613,
3.90291,
4.24711,
4.18282,
4.32505,
4.32343,
4.20834,
4.15048,
4.65123,
4.11855,
4.12835,
4.30041,
4.87421,
4.5542,
4.77747,
3.53164,
4.54348,
3.97912,
4.61723,
4.20526,
3.86804,
4.58513,
2.4436,
4.49121,
4.57528,
4.8978,
1.81068,
3.86554,
4.74381,
2.07213,
2.09223,
3.97211,
4.83585,
4.01325,
4.81149,
4.29262,
3.87846,
4.5924,
4.15907,
4.80563,
4.26264,
4.66798,
4.2186,
4.58156,
4.75406,
3.91867,
3.60931,
3.50607,
4.30856,
4.55824,
4.73856,
3.77214,
4.7273,
4.50153,
4.54082,
3.99183,
4.69438,
4.25034,
4.32047,
3.75278,
4.90787,
4.97139,
3.96534,
4.03482,
4.74396,
4.56518,
4.30262,
4.01339,
4.93153,
4.89096,
4.65489,
4.73062,
3.94436,
4.1008,
4.85157,
4.89386,
4.25616,
4.71778,
4.52003,
4.08321,
4.05076,
4.46609,
4.57562,
4.73654,
4.70187,
4.57039,
4.77104,
3.93438,
4.81294,
4.23231,
3.85885,
4.69757,
4.14618,
4.4767,
4.20894,
4.26666,
4.69035,
4.71914,
4.65206,
4.00772,
4.99633,
4.7842,
4.57934,
4.25921,
4.92866,
4.92066,
4.84729,
4.07633,
4.69198,
4.8472,
4.36999,
4.30751,
4.59363,
4.89443,
4.97367,
4.65698,
4.75577,
4.94081,
4.42736,
4.81546,
4.90015,
3.8865,
4.22402,
3.97673,
3.77515,
4.01886,
4.39418,
4.69483,
4.23938,
3.93408,
4.32132,
4.09313,
4.27052,
3.77581,
3.90642,
4.87223,
4.13688,
4.5701,
4.06878,
3.81606,
4.18979,
4.63066,
4.53284,
3.91224,
4.71342,
4.96212,
4.32695,
4.98233,
3.79912,
4.82097,
4.726,
3.76174,
4.78376,
4.83629,
4.48898,
4.21947,
3.99312,
3.74855,
4.15266,
3.97028,
2.44914,
4.48649,
4.4943,
4.48676,
1.80093,
3.84543,
4.14906,
3.64568,
4.20456,
2.0634,
2.08226,
3.69454,
4.70135,
4.96654,
4.13868,
4.82714,
4.69567,
4.72155,
4.00437,
4.83894,
4.34895,
4.07683,
4.85,
4.69759,
3.69614,
3.69552,
4.09989,
4.79662,
4.08742,
4.39171,
4.90438,
4.72757,
3.88204,
4.43897,
4.66711,
4.68764,
4.64031,
4.45104,
3.9801,
4.23864,
4.47312,
4.38623,
4.28261,
3.5855,
4.8045,
4.82138,
4.81575,
3.62252,
4.27848,
4.54622,
4.01775,
4.61043,
4.30651,
4.56837,
4.68532,
4.35168,
4.61023,
4.75734,
4.10411,
4.92689,
4.41373,
4.8445,
4.22523,
4.93041,
4.57219,
3.78393,
3.64814,
4.40099,
4.17141,
4.69466,
4.33419,
4.11137,
4.61878,
4.55391,
4.17407,
3.90412,
4.40764,
4.28297,
4.51421,
3.90996,
4.61575,
3.91039,
4.4485,
4.43099,
4.51967,
3.72261,
4.46829,
4.38155,
4.84554,
4.22733,
4.25335,
4.35288,
4.86008,
4.393,
4.9573,
4.42847,
3.99291,
4.75275,
3.89117,
4.49308,
4.84515,
4.53351,
4.94761,
4.02777,
4.75923,
4.8057,
4.77007,
3.84847,
4.24137,
4.6375,
4.57668,
4.47105,
4.26042,
4.44931,
4.25197,
3.89163,
4.04561,
4.82765,
4.61711,
4.59457,
4.61138,
4.98904,
4.95279,
4.21255,
4.76795,
4.77212,
4.77864,
4.2553,
4.29399,
4.79407,
4.68346,
4.00452,
4.61783,
4.77926,
4.8671,
3.77992,
4.67671,
4.81343,
4.98756,
3.83993,
4.58625,
4.56616,
4.3201,
4.19796,
4.20056,
4.98556,
4.40154,
4.80278,
4.00618,
4.30136,
4.46186,
4.76943,
3.69099,
4.5102,
4.37422,
3.83429,
4.55511,
3.74574,
4.69465,
4.43827,
4.99173,
3.96379,
4.54558,
4.0102,
4.45755,
2.45303,
4.49611,
4.07024,
1.80418,
3.8829,
4.50008,
2.09761,
2.09195,
4.1892,
3.40327,
4.53171,
4.99973,
3.95114,
4.34065,
3.97661,
4.90314,
4.91379,
4.47745,
4.49318,
4.56029,
4.22966,
4.29272,
4.37822,
4.43362,
4.73683,
3.94762,
4.2354,
2.96942,
3.06796,
2.08936,
4.91172,
4.66984,
3.07717,
4.35063,
4.11422,
3.44146,
4.62576,
4.81553,
4.7342,
3.71716,
4.09466,
4.55791,
4.07394,
4.86948,
4.21349,
4.60791,
4.40358,
4.74247,
4.94861,
4.1499,
4.48254,
4.63105,
4.23025,
4.20469,
4.21,
4.54222,
3.95919,
3.70554,
4.34998,
4.37754,
4.95452,
4.56624,
4.85811;
}
