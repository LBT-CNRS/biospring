netcdf SpringNetwork {

dimensions:
	spatialdim = 3;
	particle_number = 2586;
	particlename_length = 5;
	chainname_length = 4;
	resname_length = 4;

variables:
	float   coordinates(particle_number, spatialdim); 
	        coordinates:units = "angstrom" ;
	        coordinates:long_name = "Particle coordinates";

	int     particleids(particle_number); 
	        particleids:long_name = "Particle ids in source database";

	char    particlenames(particle_number,particlename_length); 
	        particlenames:long_name = "Particle name";

	float   charges(particle_number);
	        charges:long_name = "Particle charge id";
	        charges:units = "electron" ;

	float   radii(particle_number);
	        radii:units = "A" ;
	        radii:long_name = "Particle radius";

	float   epsilon(particle_number);
	        epsilon:units = "kJ.mol-1" ;
	        epsilon:long_name = "Particle epsilon for Lennard-Jones";

	float   mass(particle_number);
	        mass:units = "Da" ;
	        mass:long_name = "Particle mass";

	float   surfaceaccessibility(particle_number);
	        surfaceaccessibility:units = "A2 or percent" ;
	        surfaceaccessibility:long_name = "Particle surface accessibility";

	float   hydrophobicityscale(particle_number);
	        hydrophobicityscale:units = "kJ.mol-1" ;
	        hydrophobicityscale:long_name = "Particle hydrophobicity scale (transfer energy)";

	char    resnames(particle_number,resname_length); 
	        resnames:long_name = "particle residue name";

	int     resids(particle_number); 
	        resids:long_name = "particle residue id";

	char    chainnames(particle_number,chainname_length); 
	        chainnames:long_name = "Chain name ";

	byte    dynamicstate(particle_number); 
	        dynamicstate:long_name = "particle dynamic state (static 0 or dynamic 1)";

	int     nbspringsperparticle(particle_number); 
	        nbspringsperparticle:long_name = "Number of springs per particle";

data:
	particleids = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	coordinates = 
-2.647, -6.526, -17.499,
-1.836, -6.727, -16.646,
-2.251, -5.272, -18.209,
-1.601, -5.618, -19.15,
-3.44, -4.507, -18.793,
-3.76, -4.204, -17.685,
-4.581, -4.482, -19.154,
-3.135, -3.808, -20.104,
-3.623, -4.302, -21.077,
-1.988, -3.712, -20.421,
-3.665, -2.09, -20.185,
-2.831, -1.587, -21.723,
-3.257, -2.433, -22.434,
-1.827, -1.421, -21.036,
-2.763, -0.773, -22.603,
-1.46, -4.344, -17.297,
-1.916, -3.252, -16.972,
-0.212, -4.707, -17.012,
0.325, -5.479, -17.741,
0.62, -3.868, -16.162,
-0.071, -4.006, -15.202,
1.844, -4.617, -15.672,
2.103, -5.417, -16.523,
2.829, -3.961, -15.538,
1.707, -5.277, -14.683,
1.024, -2.617, -16.931,
0.963, -2.531, -18.151,
1.463, -1.621, -16.185,
1.586, -1.601, -14.708,
2.496, -1.936, -14.017,
0.717, -2.187, -14.133,
1.701, -0.105, -14.476,
0.551, 0.135, -14.284,
2.155, 0.23, -13.426,
2.448, 0.428, -15.675,
3.585, 0.585, -16,
2.242, 1.598, -15.525,
1.921, -0.392, -16.837,
0.979, 0.05, -17.414,
2.985, -0.759, -17.874,
3.655, -1.784, -17.741,
3.16, 0.023, -18.928,
2.291, 0.822, -19.059,
4.125, -0.12, -19.975,
3.929, -1.234, -20.354,
3.958, 0.97, -21.066,
4.97, 1.28, -21.623,
3.372, 1.954, -20.738,
3.017, 0.425, -22.16,
3.551, -0.477, -22.743,
2.013, -0.085, -21.755,
2.748, 1.46, -23.232,
2.993, 2.621, -23.089,
3.485, 1.192, -24.14,
1.383, 1.292, -23.87,
1.411, 1.585, -25.033,
0.943, 0.18, -23.945,
0.316, 2.166, -23.305,
0.655, 3.075, -22.607,
-0.451, 1.512, -22.663,
-0.347, 2.715, -24.141,
5.557, -0.06, -19.443,
5.831, 0.602, -18.442,
6.481, -0.7, -20.154,
6.256, -1.075, -21.26,
7.838, -0.8, -19.765,
7.679, -1.54, -18.845,
8.751, -1.542, -20.746,
9.937, -1.525, -20.609,
8.608, -1.178, -21.877,
8.52, -3.033, -20.75,
7.567, -3.557, -20.152,
9.335, -3.715, -21.406,
8.548, 0.332, -19.138,
8.959, -0.007, -17.945,
8.937, 1.509, -19.524,
8.788, 1.88, -20.644,
9.75, 2.248, -18.465,
10.08, 1.817, -17.407,
11.145, 2.548, -18.972,
11.017, 2.954, -20.092,
11.983, 3.325, -18.618,
11.92, 1.219, -19.094,
11.827, 0.542, -20.133,
12.626, 0.845, -18.029,
13.371, 0.104, -18.605,
13.16, 0.724, -16.971,
8.976, 3.434, -17.987,
9.441, 4.579, -18.083,
7.762, 3.132, -17.478,
7.453, 2.079, -17.036,
6.844, 4.173, -17.038,
7.4, 5.214, -17.209,
5.552, 4.093, -17.88,
4.586, 4.66, -17.477,
5.876, 4.395, -19.36,
5.752, 3.736, -20.351,
5.317, 5.433, -19.533,
6.997, 4.78, -19.555,
5.026, 2.779, -17.841,
4.366, 2.627, -18.805,
6.489, 4.193, -15.566,
6.677, 3.284, -14.768,
5.944, 5.327, -15.172,
5.697, 6.208, -15.93,
5.511, 5.661, -13.86,
6.082, 4.971, -13.089,
5.929, 7.1, -13.49,
5.652, 7.603, -12.443,
5.66, 7.999, -14.232,
7.414, 7.261, -13.612,
8.145, 7.506, -14.745,
7.914, 8.177, -15.699,
9.478, 7.567, -14.415,
10.314, 8.061, -15.1,
9.63, 7.361, -13.071,
10.776, 7.334, -12.282,
11.849, 7.698, -12.641,
10.606, 7.101, -10.937,
11.53, 7.241, -10.202,
9.331, 6.886, -10.375,
9.33, 6.917, -9.187,
8.204, 6.911, -11.16,
7.366, 7.448, -10.511,
8.346, 7.161, -12.527,
3.988, 5.62, -13.704,
3.287, 5.775, -14.693,
3.599, 5.481, -12.426,
4.337, 5.645, -11.517,
2.187, 5.549, -12.083,
1.75, 6.458, -12.711,
1.55, 4.192, -12.233,
0.414, 4.032, -11.916,
1.729, 3.832, -13.352,
2.179, 3.104, -11.381,
3.277, 2.395, -11.891,
3.898, 2.632, -12.872,
3.841, 1.37, -11.158,
4.639, 0.659, -11.665,
3.358, 1.059, -9.908,
3.97, 0.044, -9.212,
5.127, 0.086, -9.452,
2.277, 1.753, -9.372,
2.317, 1.898, -8.198,
1.696, 2.754, -10.113,
0.928, 3.435, -9.524,
2.054, 6.129, -10.667,
3.038, 6.18, -9.914,
0.864, 6.567, -10.305,
0.109, 7.084, -11.057,
0.531, 7.071, -8.994,
1.116, 6.457, -8.169,
0.49, 8.609, -8.775,
-0.023, 9.201, -7.871,
1.846, 9.225, -8.847,
2.308, 9.19, -7.738,
1.792, 10.422, -8.966,
2.791, 8.963, -9.532,
-0.373, 9.207, -9.762,
0.219, 10.051, -10.337,
-0.91, 6.606, -8.669,
-1.716, 6.407, -9.564,
-1.22, 6.556, -7.394,
-0.836, 7.442, -6.7,
-2.54, 6.228, -6.94,
-3.208, 7.094, -7.426,
-2.698, 5.055, -6.909,
-2.819, 6.586, -5.489,
-1.983, 7.04, -4.717,
-4.058, 6.262, -5.098,
-4.977, 6.43, -5.832,
-4.52, 6.537, -3.74,
-3.73, 6.796, -2.9,
-5.305, 7.888, -3.803,
-5.468, 8.488, -2.777,
-6.434, 7.747, -4.18,
-4.876, 8.772, -4.491,
-5.333, 5.358, -3.287,
-5.794, 4.545, -4.1,
-5.536, 5.188, -1.994,
-5.709, 6.208, -1.41,
-6.319, 4.04, -1.517,
-7.258, 4.207, -2.232,
-5.439, 2.824, -1.277,
-4.99, 2.468, -2.323,
-6.152, 1.937, -0.933,
-4.196, 3.052, -0.4,
-3.492, 3.915, -0.823,
-4.653, 3.35, 0.66,
-3.366, 1.765, -0.229,
-2.519, 1.813, -1.075,
-3.927, 0.778, -0.595,
-2.599, 1.676, 1.044,
-3.329, 1.918, 1.952,
-1.806, 2.554, 0.88,
-1.728, 0.483, 1.307,
-1.164, 0.504, 2.355,
-0.879, 0.542, 0.464,
-2.216, -0.591, 1.14,
-7.054, 4.442, -0.246,
-6.7, 5.378, 0.442,
-8.108, 3.734, 0.05,
-8.837, 3.357, -0.807,
-8.861, 3.843, 1.279,
-8.595, 4.652, 2.103,
-10.348, 4.116, 1.014,
-10.926, 4.101, 2.064,
-10.982, 3.287, 0.429,
-10.544, 5.437, 0.243,
-10.09, 5.602, -0.848,
-11.972, 5.705, -0.117,
-12.773, 5, 0.428,
-12.201, 5.592, -1.29,
-12.461, 6.782, 0.096,
-9.953, 6.529, 1.144,
-10.256, 6.461, 2.301,
-10.533, 7.563, 0.93,
-8.875, 6.89, 0.777,
-8.656, 2.483, 1.973,
-8.857, 1.403, 1.386,
-8.254, 2.519, 3.237,
-7.207, 3.059, 3.391,
-8.046, 1.237, 3.906,
-7.643, 0.519, 3.05,
-7.054, 1.308, 4.576,
-8.877, 1.072, 5.157,
-9.37, 2.041, 5.701,
-9.024, -0.162, 5.577,
-9.172, -1.054, 4.815,
-9.682, -0.552, 6.777,
-9.348, 0.381, 7.426,
-11.144, -0.927, 6.743,
-11.35, -1.175, 7.895,
-12.185, -0.422, 6.436,
-11.526, -2.155, 6.007,
-11.662, -3.422, 6.5,
-11.608, -3.874, 7.596,
-12.034, -4.308, 5.527,
-12.72, -5.209, 5.892,
-12.135, -3.614, 4.342,
-12.466, -4.071, 3.062,
-13.305, -4.911, 2.983,
-12.487, -3.149, 2.047,
-13.099, -3.449, 1.073,
-12.199, -1.782, 2.288,
-12.495, -0.904, 1.549,
-11.873, -1.345, 3.55,
-11.978, -0.17, 3.687,
-11.834, -2.265, 4.605,
-8.859, -1.671, 7.445,
-8.336, -2.595, 6.857,
-8.749, -1.512, 8.75,
-8.328, -0.484, 9.155,
-8.073, -2.521, 9.551,
-8.071, -3.523, 8.907,
-6.699, -2.081, 10.005,
-6.552, -1.399, 10.964,
-6.091, -1.637, 9.081,
-6.049, -3.222, 10.514,
-5.45, -3.677, 9.617,
-8.959, -2.837, 10.754,
-9.314, -1.915, 11.484,
-9.288, -4.099, 10.922,
-8.981, -4.978, 10.181,
-10.143, -4.582, 11.983,
-10.981, -3.742, 12.046,
-10.607, -6.018, 11.631,
-9.811, -6.882, 11.855,
-10.928, -6.257, 10.502,
-11.763, -6.486, 12.486,
-11.806, -6.668, 13.665,
-12.086, -7.554, 12.046,
-13.038, -5.702, 12.296,
-14.094, -6.166, 12.748,
-13.012, -4.543, 11.65,
-14.154, -4.193, 11.686,
-12.805, -4.536, 10.475,
-9.631, -4.569, 13.399,
-10.391, -4.809, 14.362,
-8.386, -4.352, 13.666,
-7.694, -4.356, 12.703,
-7.679, -4.27, 14.922,
-8.272, -3.315, 15.305,
-8.047, -5.279, 16.001,
-7.268, -5.024, 16.87,
-9.046, -5.424, 16.643,
-7.916, -6.729, 15.583,
-6.664, -7.305, 15.424,
-5.772, -7.096, 16.181,
-6.511, -8.61, 15.009,
-5.593, -9.274, 15.371,
-7.636, -9.371, 14.76,
-7.505, -10.682, 14.355,
-6.657, -10.739, 13.535,
-8.897, -8.832, 14.913,
-9.778, -9.602, 14.699,
-9.029, -7.517, 15.323,
-10.103, -7.518, 15.836,
-6.209, -4.33, 14.47,
-5.832, -5.241, 13.72,
-5.427, -3.305, 14.775,
-6.048, -2.959, 15.725,
-4.024, -3.326, 14.313,
-3.725, -4.369, 13.832,
-3.659, -2.048, 13.602,
-2.732, -1.566, 14.186,
-4.293, -1.127, 13.204,
-3.101, -2.168, 12.224,
-3.69, -2.889, 11.213,
-4.043, -3.993, 11.454,
-2.967, -2.789, 10.113,
-2.632, -3.167, 9.04,
-1.915, -2.04, 10.368,
-1.976, -1.633, 11.679,
-1.049, -0.97, 12.011,
-3.138, -3.585, 15.531,
-1.923, -3.667, 15.46,
-3.819, -3.716, 16.664,
-4.598, -2.92, 17.058,
-3.22, -3.952, 17.96,
-2.392, -4.808, 17.962,
-2.728, -2.624, 18.548,
-1.98, -2.578, 19.482,
-1.977, -2.128, 17.758,
-3.788, -1.578, 18.799,
-4.936, -1.901, 19.185,
-3.487, -0.372, 18.627,
-4.215, -4.615, 18.912,
-5.016, -5.48, 18.561,
-4.194, -4.205, 20.154,
-3.08, -4.12, 20.568,
-4.919, -4.485, 21.331,
-5.4, -3.4, 21.446,
-6.022, -5.539, 21.347,
-6.357, -6.014, 22.391,
-7.302, -5.048, 20.681,
-7.357, -4.293, 19.76,
-8.037, -4.568, 21.496,
-7.893, -6.033, 20.336,
-5.611, -6.773, 20.759,
-4.563, -7.082, 21.219,
-3.95, -4.807, 22.5,
-3.41, -3.87, 23.091,
-5.121, -3.794, 23.764,
-6.203, -3.345, 23.579,
-4.737, -3.232, 25.134,
-3.583, -2.913, 25.153,
-5.211, -2.141, 25.255,
-4.643, -4.176, 26.396,
-3.543, -4.775, 26.542,
-5.768, -4.019, 27.193,
-6.262, -2.941, 27.122,
-6.353, -4.742, 28.463,
-7.234, -3.961, 28.639,
-6.547, -6.228, 28.185,
-5.465, -6.711, 28.016,
-6.962, -6.852, 29.115,
-7.389, -6.485, 26.922,
-6.811, -6.212, 25.916,
-7.646, -7.972, 26.658,
-8.292, -8.57, 27.472,
-6.643, -8.629, 26.593,
-8.172, -8.233, 25.612,
-8.778, -5.834, 26.958,
-9.158, -5.736, 28.082,
-8.81, -4.842, 26.29,
-9.648, -6.476, 26.438,
-5.647, -4.652, 29.913,
-4.417, -4.528, 30.019,
-6.587, -4.757, 30.984,
-7.708, -4.462, 30.745,
-6.359, -4.832, 32.54,
-5.248, -5.267, 32.583,
-6.704, -3.506, 33.216,
-7.788, -3.05, 33.03,
-6.491, -3.544, 34.736,
-6.284, -4.588, 35.284,
-5.559, -2.936, 35.189,
-7.417, -3.087, 35.345,
-5.834, -2.349, 32.711,
-5.56, -1.775, 31.689,
-4.761, -2.89, 32.768,
-6.106, -1.03, 33.433,
-6.392, -0.135, 32.684,
-7.007, -0.872, 34.207,
-5.142, -0.606, 34.009,
-7.167, -5.984, 33.05,
-8.337, -6.17, 32.676,
-6.687, -6.866, 33.965,
-5.631, -7.107, 34.46,
-7.581, -7.959, 33.931,
-7.103, -8.922, 33.41,
-8.385, -8.259, 35.186,
-9.117, -7.878, 36.049,
-9.048, -9.19, 34.819,
-7.646, -9.041, 36.268,
-6.907, -9.97, 35.96,
-7.82, -8.72, 37.538,
-6.816, -8.69, 38.18,
-8.718, -8.888, 38.302,
-8.633, -7.35, 33.071,
-8.496, -7.38, 31.826,
-9.436, -6.789, 33.941,
-8.887, -6.054, 34.702,
-10.626, -5.981, 33.749,
-11.503, -6.777, 33.905,
-10.721, -5.053, 34.976,
-11.234, -4.239, 34.254,
-11.034, -4.216, 35.79,
-10.564, -5.814, 36.315,
-11.419, -6.637, 36.654,
-9.525, -5.597, 37.107,
-8.4, -5.244, 37.265,
-9.966, -5.435, 38.207,
-10.558, -5.188, 32.446,
-9.647, -4.374, 32.239,
-11.567, -5.467, 31.636,
-12.575, -5.867, 32.125,
-11.749, -4.905, 30.279,
-10.78, -5.323, 29.736,
-12.969, -5.575, 29.648,
-14.015, -5.248, 30.127,
-13.112, -5.39, 28.477,
-12.851, -7.104, 29.675,
-11.893, -7.654, 29.131,
-13.767, -7.832, 30.284,
-14.365, -7.833, 31.313,
-14.197, -8.744, 29.647,
-11.91, -3.368, 30.316,
-12.432, -2.805, 31.288,
-11.446, -2.737, 29.222,
-10.845, -3.306, 28.374,
-11.435, -1.248, 29.051,
-10.316, -0.838, 29.132,
-12.005, -0.7, 29.946,
-12.27, -0.813, 27.827,
-13.372, -0.275, 27.987,
-12.009, -0.977, 26.397,
-10.54, -1.045, 26.144,
-9.968, -0.103, 26.605,
-9.889, -1.967, 26.533,
-10.456, -1.174, 24.652,
-10.343, -2.32, 24.328,
-9.487, -0.653, 24.182,
-11.724, -0.6, 24.116,
-11.74, 0.593, 24.04,
-11.764, -0.897, 22.96,
-12.782, -0.907, 25.162,
-13.653, -0.132, 25.407,
-13.535, -2.184, 24.851,
-13.382, -3.182, 25.57,
-14.363, -2.201, 23.798,
-14.497, -1.188, 23.193,
-15.133, -3.394, 23.455,
-15.088, -4.27, 24.267,
-16.647, -3.12, 23.365,
-17.358, -4.077, 23.284,
-17.149, -2.307, 24.556,
-18.344, -2.289, 24.455,
-16.88, -1.172, 24.811,
-16.998, -2.887, 25.594,
-16.985, -2.425, 22.159,
-15.999, -2.012, 21.666,
-14.65, -4.156, 22.23,
-14.869, -5.378, 22.124,
-13.996, -3.533, 21.277,
-13.093, -2.912, 21.737,
-13.456, -4.121, 20.051,
-12.517, -4.778, 20.384,
-14.458, -4.967, 19.312,
-15.46, -4.321, 19.229,
-14.207, -5.164, 18.158,
-14.718, -6.355, 19.672,
-15.837, -6.545, 20.145,
-17.008, -6.345, 20.226,
-15.62, -7.848, 20.427,
-16.283, -8.704, 20.917,
-14.403, -8.217, 20.017,
-13.784, -7.101, 19.424,
-12.857, -7.56, 18.838,
-12.934, -2.97, 19.193,
-13.127, -1.826, 19.673,
-12.291, -3.152, 18.031,
-11.876, -4.197, 17.647,
-11.822, -1.904, 17.388,
-12.853, -1.306, 17.469,
-10.543, -1.421, 18.035,
-10.54, -1.678, 19.204,
-10.686, -0.238, 18.079,
-9.2, -1.87, 17.514,
-9.111, -1.515, 16.386,
-9.161, -2.997, 17.901,
-8.072, -1.206, 18.304,
-8.17, -1.131, 19.551,
-7.087, -0.741, 17.704,
-11.762, -1.868, 15.885,
-11.698, -2.834, 15.155,
-11.842, -0.639, 15.354,
-12.146, 0.325, 15.977,
-11.834, -0.406, 13.93,
-11.613, -1.391, 13.305,
-13.23, -0.065, 13.393,
-13.853, 0.803, 13.924,
-13.261, 0.235, 12.235,
-14.144, -1.264, 13.268,
-13.877, -2.155, 12.447,
-15.2, -1.265, 14.082,
-15.544, -0.791, 15.116,
-16.121, -1.926, 13.713,
-10.945, 0.794, 13.591,
-11.058, 1.824, 14.247,
-10.124, 0.604, 12.569,
-9.694, -0.49, 12.673,
-9.279, 1.638, 12.034,
-9.829, 2.592, 12.48,
-7.789, 1.39, 12.121,
-7.373, 0.733, 11.224,
-7.48, 2.516, 11.855,
-7.163, 1.298, 13.481,
-6.107, 1.809, 13.259,
-7.736, 1.812, 14.387,
-6.888, -0.173, 13.805,
-6.313, -0.791, 12.972,
-7.937, -0.703, 13.991,
-6.044, -0.313, 15.054,
-5.225, -1.093, 15.413,
-6.911, -0.141, 15.852,
-5.218, 0.892, 15.338,
-4.565, 0.646, 16.315,
-4.384, 1.044, 14.495,
-5.759, 1.873, 15.75,
-9.606, 1.791, 10.527,
-9.752, 0.806, 9.826,
-9.663, 3.019, 10.094,
-9.991, 3.928, 10.784,
-9.909, 3.417, 8.748,
-9.456, 2.509, 8.137,
-11.251, 4.197, 8.592,
-11.389, 5.11, 9.354,
-11.35, 4.793, 7.559,
-12.45, 3.235, 8.717,
-12.62, 2.592, 9.707,
-13.726, 3.997, 8.592,
-13.806, 5.048, 8.016,
-14.225, 4.226, 9.656,
-14.615, 3.386, 8.064,
-12.351, 2.207, 7.586,
-12.592, 2.623, 6.487,
-13.253, 1.44, 7.776,
-11.369, 1.557, 7.514,
-8.834, 4.424, 8.353,
-8.431, 5.191, 9.213,
-8.45, 4.408, 7.079,
-8.431, 3.607, 6.216,
-7.491, 5.389, 6.645,
-8.067, 6.416, 6.863,
-6.402, 5.117, 7.012,
-7.381, 5.442, 5.128,
-8.136, 4.898, 4.348,
-6.306, 6.109, 4.749,
-5.77, 6.857, 5.496,
-6.017, 6.36, 3.367,
-6.282, 5.384, 2.749,
-6.606, 7.762, 3.132,
-6.446, 8.42, 2.142,
-6.37, 8.533, 4.01,
-7.801, 7.719, 3.201,
-4.53, 6.322, 3.131,
-3.771, 6.127, 4.088,
-4.117, 6.478, 1.879,
-4.746, 7.238, 1.218,
-2.686, 6.398, 1.563,
-2.341, 5.261, 1.56,
-2.279, 7.362, 2.134,
-2.491, 6.795, 0.116,
-3.476, 6.907, -0.6,
-1.255, 7.052, -0.275,
-0.559, 7.685, 0.447,
-0.955, 7.453, -1.642,
-1.827, 7.203, -2.398,
-0.654, 8.949, -1.767,
-1.266, 9.505, -2.637,
0.468, 9.316, -1.977,
-0.963, 9.639, -0.836,
0.263, 6.631, -2.051,
1.041, 6.277, -1.146,
0.399, 6.319, -3.333,
0.311, 7.342, -3.933,
1.578, 5.52, -3.679,
2.396, 6.166, -3.105,
1.321, 3.979, -3.588,
2.223, 3.238, -3.825,
1.019, 3.73, -2.462,
0.162, 3.521, -4.429,
-1.139, 3.52, -3.917,
-1.365, 3.581, -2.756,
-2.187, 3.114, -4.75,
-3.275, 3.062, -4.287,
-1.962, 2.725, -6.062,
-2.955, 2.238, -6.487,
-0.671, 2.719, -6.579,
-0.549, 2.56, -7.743,
0.387, 3.13, -5.749,
1.453, 3.209, -6.257,
2.006, 5.918, -5.085,
1.167, 6.392, -5.851,
3.275, 5.691, -5.374,
4.01, 6.302, -4.666,
3.747, 6.006, -6.758,
4.437, 6.969, -6.57,
3.153, 6.298, -7.738,
4.766, 4.889, -7.067,
5.345, 4.309, -6.135,
4.93, 4.594, -8.355,
5.278, 5.628, -8.832,
5.866, 3.533, -8.704,
5.244, 2.529, -8.608,
6.829, 3.902, -8.099,
6.434, 3.679, -10.089,
6.112, 4.532, -10.913,
7.356, 2.788, -10.386,
8.179, 2.559, -9.563,
8.026, 2.699, -11.672,
7.493, 3.365, -12.493,
9.447, 3.207, -11.571,
10.165, 2.789, -10.711,
9.472, 4.364, -11.283,
10.273, 3.072, -12.811,
10.09, 3.93, -13.902,
9.527, 4.967, -13.86,
10.869, 3.81, -15.031,
11.163, 4.794, -15.631,
11.837, 2.83, -15.102,
12.61, 2.703, -16.237,
13.545, 3.418, -16.083,
12.044, 1.972, -14.047,
13.175, 1.624, -13.912,
11.262, 2.094, -12.907,
11.912, 1.766, -11.967,
7.943, 1.242, -12.121,
8.256, 0.344, -11.354,
7.45, 1.042, -13.334,
8, 1.719, -14.137,
7.365, -0.32, -13.878,
7.036, -0.982, -12.948,
6.121, -0.439, -14.752,
5.287, 0.219, -14.208,
6.423, 0.161, -15.737,
5.584, -1.835, -14.93,
5.961, -2.882, -15.373,
5.197, -1.557, -16.028,
5.031, -2.515, -13.726,
4.357, -1.94, -12.881,
5.299, -3.819, -13.617,
4.602, -4.725, -13.947,
5.629, -4.165, -12.529,
8.647, -0.643, -14.637,
9.152, 0.202, -15.386,
9.232, -1.807, -14.444,
9.344, -1.9, -13.27,
10.48, -2.134, -15.172,
11.059, -1.216, -15.662,
11.511, -2.86, -14.287,
11.16, -3.922, -13.897,
12.722, -3.293, -15.099,
13.528, -3.873, -14.423,
12.673, -3.997, -16.067,
13.391, -2.383, -15.508,
11.954, -1.922, -13.149,
13.089, -1.555, -13.295,
12.05, -2.591, -12.163,
11.423, -0.897, -12.846,
10.149, -2.968, -16.412,
10.665, -2.732, -17.496,
9.276, -3.928, -16.256,
9.208, -4.377, -15.166,
8.782, -4.822, -17.297,
8.417, -4.091, -18.157,
9.807, -5.869, -17.622,
10.711, -5.265, -18.125,
9.887, -6.785, -18.39,
10.1, -6.782, -16.428,
9.202, -7.355, -15.817,
11.365, -6.935, -16.055,
12.315, -6.436, -15.544,
11.81, -7.997, -16.375,
7.447, -5.338, -16.785,
7.055, -5.019, -15.665,
6.703, -6.14, -17.504,
7.015, -6.562, -18.905,
7.972, -7.055, -19.427,
6.715, -5.686, -19.663,
5.93, -7.57, -19.221,
6.339, -8.693, -19.17,
5.687, -7.491, -20.393,
4.8, -7.349, -18.288,
3.703, -7.12, -17.856,
4.229, -8.153, -18.98,
5.378, -6.559, -17.103,
4.841, -5.495, -17.11,
5.289, -7.316, -15.825,
4.178, -7.545, -15.31,
6.362, -7.803, -15.278,
7.114, -8.159, -16.121,
6.321, -8.615, -14.075,
5.229, -9.008, -13.819,
7.247, -9.837, -14.342,
8.423, -9.856, -14.558,
7.227, -10.618, -13.433,
6.75, -10.585, -15.558,
5.642, -11.412, -15.43,
5.517, -12.107, -14.474,
5.144, -12.104, -16.512,
4.796, -13.24, -16.483,
5.761, -11.958, -17.755,
5.219, -12.659, -18.824,
6.018, -12.712, -19.694,
6.845, -11.126, -17.903,
7.521, -11.226, -18.877,
7.343, -10.431, -16.804,
8.52, -10.389, -16.979,
6.819, -7.876, -12.85,
6.458, -8.322, -11.76,
7.671, -6.84, -13.019,
8.076, -6.371, -14.023,
8.274, -6.172, -11.919,
7.502, -6.466, -11.067,
9.686, -6.707, -11.565,
9.743, -6.984, -10.406,
10.175, -7.912, -12.333,
10.065, -8.932, -11.712,
9.842, -8.25, -13.427,
11.371, -7.971, -12.46,
10.776, -5.666, -11.615,
10.643, -4.619, -11.055,
11.405, -5.681, -12.63,
11.661, -6.099, -10.921,
8.254, -4.644, -11.976,
8.555, -3.965, -12.957,
7.897, -4.086, -10.807,
7.914, -4.683, -9.789,
7.821, -2.648, -10.555,
8.638, -2.049, -11.169,
6.654, -2.421, -10.495,
8.309, -2.377, -9.127,
8.517, -3.274, -8.287,
8.584, -1.126, -8.838,
9.157, -0.432, -9.609,
9.008, -0.721, -7.494,
8.748, -1.589, -6.731,
10.444, -0.198, -7.507,
10.687, 0.765, -8.174,
10.872, 0.187, -6.458,
11.371, -1.333, -7.848,
11.58, -2.342, -6.948,
11.994, -1.949, -5.901,
12.432, -3.397, -7.236,
13.139, -3.957, -6.46,
13.055, -3.41, -8.476,
13.907, -4.215, -8.682,
12.833, -2.404, -9.391,
13.841, -2.204, -9.992,
11.981, -1.363, -9.089,
12.415, -0.361, -9.563,
8.096, 0.418, -7.045,
7.838, 1.301, -7.87,
7.598, 0.42, -5.821,
8.462, 0.266, -5.024,
6.756, 1.531, -5.42,
7.352, 2.393, -5.988,
5.24, 1.317, -5.439,
4.795, 1.971, -6.328,
4.711, 1.615, -4.41,
4.728, -0.049, -5.616,
5.194, -0.625, -6.551,
4.927, -0.747, -4.672,
3.219, -0.103, -5.813,
2.537, 0.123, -4.78,
2.711, -0.387, -6.929,
7.075, 1.997, -3.995,
7.551, 1.382, -3.062,
6.633, 3.217, -3.882,
6.819, 3.981, -4.77,
6.717, 4, -2.685,
7.389, 3.483, -1.859,
7.529, 5.252, -3.133,
7.1, 6.032, -3.932,
8.652, 5.057, -3.506,
7.893, 6.085, -1.922,
7.746, 7.233, -2.225,
7.525, 5.978, -0.798,
9.666, 6.276, -1.731,
9.693, 7.131, -0.128,
10.864, 6.905, -0.046,
9.574, 8.283, -0.418,
9.218, 6.93, 0.944,
5.312, 4.394, -2.275,
4.53, 4.881, -3.091,
4.982, 4.221, -0.999,
5.824, 4.334, -0.179,
3.711, 4.676, -0.511,
3.038, 3.692, -0.502,
3.593, 5.665, -1.161,
3.773, 5.275, 0.888,
4.641, 5.006, 1.699,
2.729, 6.049, 1.167,
2.615, 6.908, 0.355,
2.531, 6.647, 2.485,
3.376, 6.348, 3.254,
2.684, 8.185, 2.349,
3.813, 8.557, 2.203,
2.151, 8.826, 1.492,
2.185, 8.863, 3.615,
2.877, 8.744, 4.812,
3.898, 9.332, 4.632,
2.379, 9.343, 5.955,
3.174, 9.781, 6.724,
1.198, 10.06, 5.901,
0.714, 10.65, 7.042,
0.98, 11.806, 6.959,
0.486, 10.186, 4.726,
0.037, 11.279, 4.58,
0.994, 9.579, 3.585,
0.598, 10.164, 2.628,
1.14, 6.226, 2.928,
0.202, 6.334, 2.112,
0.934, 5.719, 4.112,
1.615, 6.037, 5.024,
-0.395, 5.33, 4.556,
-1.26, 5.586, 3.788,
-0.568, 3.847, 4.756,
0.198, 3.503, 5.607,
-1.643, 3.506, 5.152,
-0.313, 2.87, 3.674,
-0.453, 3.149, 2.473,
0.029, 1.716, 4.035,
-0.668, 5.961, 5.938,
0.237, 6.225, 6.727,
-1.944, 6.086, 6.247,
-2.51, 6.8, 5.491,
-2.367, 6.615, 7.542,
-1.598, 5.964, 8.173,
-2.482, 8.108, 7.561,
-2.332, 8.414, 8.7,
-1.598, 8.656, 6.976,
-3.695, 8.784, 7.095,
-4.88, 8.829, 7.782,
-5.387, 8.621, 8.835,
-5.817, 9.529, 7.055,
-6.86, 9.932, 7.461,
-5.235, 9.963, 5.886,
-5.768, 10.713, 4.84,
-6.754, 11.353, 5.02,
-4.967, 11, 3.76,
-5.371, 11.83, 3.009,
-3.638, 10.546, 3.718,
-3.048, 11.036, 2.81,
-3.115, 9.805, 4.774,
-2.019, 9.456, 4.496,
-3.912, 9.513, 5.874,
-3.619, 5.877, 7.985,
-4.473, 5.568, 7.139,
-3.674, 5.563, 9.272,
-2.842, 5.569, 10.106,
-4.8, 4.882, 9.864,
-5.724, 5.248, 9.219,
-4.484, 3.435, 10.222,
-5.134, 3.107, 11.165,
-3.367, 3.394, 10.643,
-4.465, 2.4, 9.127,
-3.687, 2.697, 8.272,
-3.925, 1.083, 9.687,
-4.719, 0.285, 10.069,
-3.229, 0.613, 8.831,
-3.129, 1.172, 10.578,
-5.855, 2.171, 8.495,
-6.296, 3.18, 8.053,
-5.641, 1.547, 7.499,
-6.697, 1.621, 9.126,
-5.201, 5.61, 11.16,
-4.344, 6.014, 11.94,
-6.476, 5.761, 11.397,
-7.15, 6.338, 10.603,
-6.996, 6.412, 12.592,
-7.702, 7.369, 12.423,
-6.199, 6.978, 13.271,
-7.978, 5.476, 13.286,
-8.735, 4.807, 12.598,
-7.941, 5.404, 14.61,
-7.968, 6.512, 15.043,
-8.913, 4.527, 15.317,
-9.059, 3.464, 14.817,
-8.496, 4.298, 16.745,
-7.968, 5.333, 17.015,
-7.761, 3.364, 16.762,
-9.56, 4.198, 17.808,
-10.731, 4.413, 17.686,
-9.423, 5.158, 18.512,
-9.716, 2.807, 18.389,
-10.21, 2.089, 17.576,
-10.524, 2.836, 19.275,
-8.608, 2.316, 19.153,
-8.106, 1.42, 18.563,
-7.837, 2.853, 20.083,
-7.964, 4.099, 20.524,
-7.16, 4.448, 21.327,
-9.073, 4.49, 20.715,
-6.869, 2.076, 20.595,
-6.56, 0.949, 20.376,
-6.181, 2.337, 21.533,
-10.273, 5.208, 15.215,
-10.317, 6.436, 15.275,
-11.325, 4.447, 14.996,
-11.483, 3.392, 15.514,
-12.672, 5.036, 14.876,
-12.404, 6.105, 14.433,
-13.484, 4.364, 13.781,
-12.863, 3.78, 12.946,
-14.205, 3.575, 14.315,
-14.18, 5.31, 12.838,
-14.774, 5.745, 11.888,
-15.27, 4.876, 13.11,
-13.091, 6.43, 11.93,
-14.011, 7.972, 12.131,
-15.184, 8.189, 12.055,
-13.61, 8.272, 11.043,
-13.461, 8.782, 12.816,
-13.391, 4.978, 16.224,
-13.384, 3.943, 16.896,
-13.978, 6.101, 16.619,
-13.991, 7.371, 15.839,
-14.289, 7.625, 14.716,
-12.966, 7.927, 16.114,
-14.985, 8.226, 16.583,
-14.753, 9.401, 16.631,
-16.054, 8.252, 16.043,
-14.994, 7.728, 17.983,
-14.243, 8.239, 18.763,
-16.058, 8.051, 18.426,
-14.645, 6.236, 17.889,
-13.845, 6.003, 18.743,
-15.89, 5.394, 18.08,
-16.871, 5.645, 17.379,
-15.856, 4.425, 18.996,
-14.908, 4.13, 19.649,
-16.952, 3.591, 19.366,
-17.699, 4.483, 19.633,
-17.572, 2.707, 18.247,
-17.729, 1.534, 18.415,
-17.01, 2.713, 17.193,
-19.002, 3.265, 18.124,
-19.979, 2.957, 19.057,
-20.148, 1.831, 19.399,
-21.247, 3.501, 18.94,
-22.175, 3.535, 19.677,
-21.523, 4.369, 17.902,
-22.779, 4.917, 17.775,
-22.653, 6.093, 17.71,
-20.541, 4.697, 16.998,
-20.829, 5.408, 16.089,
-19.29, 4.148, 17.1,
-18.802, 4.187, 16.016,
-16.788, 2.706, 20.598,
-16.177, 1.64, 20.524,
-17.397, 3.136, 21.701,
-17.538, 4.314, 21.817,
-17.385, 2.456, 22.981,
-16.582, 3.232, 23.41,
-18.757, 1.805, 23.278,
-18.837, 1.091, 24.232,
-18.828, 0.986, 22.407,
-19.902, 2.815, 23.3,
-20.027, 3.927, 23.726,
-19.987, 3.04, 22.129,
-21.226, 2.17, 23.708,
-21.461, 2.466, 24.843,
-21.326, 0.978, 23.719,
-22.362, 2.728, 22.808,
-22.479, 3.918, 22.793,
-22.32, 2.265, 21.709,
-23.713, 2.211, 23.224,
-24.552, 3.055, 23.074,
-23.9, 1.859, 24.355,
-24.137, 1.272, 22.608,
-16.281, 1.419, 23.131,
-15.296, 1.597, 23.854,
-18.053, 3.17, 25.045,
-18.031, 4.247, 24.533,
-18.083, 3.745, 26.381,
-19.073, 4.393, 26.551,
-17.069, 4.379, 26.417,
-18.038, 2.61, 27.421,
-18.231, 1.422, 27.094,
-17.791, 3.078, 28.605,
-17.895, 4.264, 28.624,
-17.527, 2.303, 29.807,
-18.483, 2.332, 30.522,
-17.37, 0.824, 29.489,
-17.073, 0.197, 30.467,
-18.332, 0.204, 29.136,
-16.268, 0.628, 28.621,
-15.75, 1.665, 28.403,
-16.251, 2.895, 30.339,
-15.257, 2.193, 30.561,
-16.365, 4.179, 30.447,
-17.398, 4.709, 30.724,
-15.325, 5.02, 30.934,
-15.685, 6.126, 30.657,
-15.029, 4.747, 32.414,
-15.036, 3.575, 32.643,
-13.838, 5.559, 32.942,
-14.234, 5.711, 34.08,
-12.868, 6.047, 33.497,
-14.186, 6.655, 32.562,
-16.195, 5.069, 33.34,
-17.15, 4.39, 33.085,
-16.154, 4.897, 34.531,
-16.66, 6.176, 33.29,
-13.995, 4.782, 30.269,
-13.198, 3.921, 30.653,
-13.624, 5.438, 29.191,
-14.229, 5.954, 28.306,
-12.199, 5.451, 29.228,
-11.936, 6.618, 29.19,
-11.841, 4.522, 30.408,
-10.7, 4.87, 30.568,
-11.55, 3.43, 29.991,
-12.793, 4.736, 31.62,
-12.813, 5.919, 31.335,
-11.725, 4.956, 32.156,
-12.56, 3.769, 32.793,
-11.693, 2.822, 32.687,
-13.232, 3.902, 33.892,
-11.25, 5.108, 28.078,
-10.139, 4.65, 28.37,
-11.66, 4.551, 24.96,
-12.34, 4.423, 24.001,
-10.602, 5.265, 25.654,
-11.323, 5.942, 26.318,
-9.387, 4.412, 25.985,
-9.172, 3.777, 26.976,
-8.44, 5.132, 26.11,
-9.221, 3.091, 25.294,
-10.071, 2.191, 25.395,
-8.117, 2.884, 24.568,
-7.029, 2.732, 25.027,
-8.253, 2.321, 23.531,
-10.208, 6.561, 24.945,
-10.913, 7.576, 25.093,
-9.092, 6.566, 24.211,
-8.451, 5.645, 23.831,
-8.654, 7.779, 23.532,
-9.531, 8.582, 23.407,
-7.837, 8.166, 24.311,
-8.177, 7.585, 22.1,
-8.362, 6.542, 21.472,
-7.533, 8.605, 21.539,
-7.721, 9.641, 22.09,
-6.997, 8.676, 20.203,
-8.009, 8.523, 19.585,
-6.617, 10.141, 19.891,
-7.401, 10.962, 20.279,
-5.532, 10.601, 20.086,
-6.715, 10.347, 18.712,
-5.813, 7.776, 19.841,
-4.894, 7.494, 20.6,
-5.828, 7.284, 18.596,
-6.537, 7.843, 17.824,
-4.824, 6.427, 18.022,
-3.833, 6.725, 18.604,
-5.053, 4.935, 18.221,
-6.039, 4.382, 17.867,
-5.012, 4.766, 19.403,
-3.968, 4.072, 17.625,
-3.919, 3.84, 16.238,
-4.627, 4.285, 15.397,
-2.947, 3.062, 15.654,
-2.967, 2.879, 14.486,
-1.981, 2.473, 16.455,
-0.992, 1.684, 15.901,
-0.256, 2.375, 15.301,
-1.997, 2.675, 17.829,
-1.214, 2.068, 18.486,
-2.989, 3.471, 18.405,
-3.271, 2.94, 19.431,
-4.682, 6.737, 16.527,
-5.622, 6.65, 15.748,
-3.46, 7.043, 16.146,
-2.49, 6.854, 16.796,
-3.136, 7.382, 14.756,
-4.042, 7.047, 14.068,
-3.079, 8.889, 14.672,
-2.694, 9.361, 15.702,
-4.215, 9.269, 14.663,
-2.349, 9.589, 13.586,
-1.272, 9.998, 13.906,
-2.187, 8.893, 12.637,
-3.051, 10.881, 13.144,
-4.238, 11.027, 13.218,
-2.733, 11.756, 13.902,
-2.677, 11.269, 11.728,
-3.127, 12.379, 11.609,
-1.526, 11.584, 11.683,
-3.405, 10.542, 10.644,
-4.565, 10.405, 10.913,
-3.465, 11.268, 9.691,
-2.886, 9.493, 10.446,
-1.853, 6.671, 14.362,
-0.878, 6.647, 15.113,
-1.816, 6.009, 13.195,
-2.426, 6.576, 12.357,
-0.591, 5.367, 12.746,
0.259, 5.955, 13.327,
-0.527, 3.877, 12.85,
0.387, 3.443, 13.483,
-1.554, 3.305, 13.021,
-0.214, 3.456, 11.77,
-0.265, 5.903, 11.361,
-1.132, 6.277, 10.601,
1.012, 5.974, 11.064,
1.904, 5.602, 11.746,
1.387, 6.484, 9.745,
0.757, 5.717, 9.082,
1.226, 7.93, 9.725,
0.962, 8.217, 8.599,
0.432, 8.286, 10.54,
2.3, 8.892, 10.136,
2.6, 8.994, 11.289,
3.358, 8.858, 9.582,
1.83, 10.324, 9.918,
2.546, 11.297, 10.027,
0.55, 10.479, 9.583,
-0.182, 11.214, 8.995,
0.279, 10.779, 10.709,
2.645, 5.781, 9.299,
3.333, 5.188, 10.152,
2.888, 5.693, 7.976,
2.814, 6.732, 7.409,
4.063, 4.917, 7.537,
3.927, 3.754, 7.738,
4.876, 5.498, 8.184,
4.405, 5.167, 6.078,
3.556, 5.423, 5.219,
5.72, 5.145, 5.813,
6.43, 5.656, 6.615,
6.236, 5.238, 4.469,
5.328, 5.412, 3.73,
7.18, 6.398, 4.146,
7.199, 6.779, 3.015,
6.66, 7.629, 4.888,
7.425, 8.027, 5.725,
6.703, 8.568, 4.139,
5.625, 7.759, 5.466,
8.601, 6.118, 4.529,
9.232, 7.107, 4.793,
8.969, 5.341, 5.352,
9.199, 5.758, 3.552,
6.868, 3.883, 4.142,
7.535, 3.264, 4.98,
6.516, 3.38, 2.946,
6.855, 4.22, 2.177,
7.007, 2.045, 2.537,
8.033, 1.998, 3.137,
5.867, 1.042, 2.666,
6.319, 0.034, 2.226,
5.533, 1.019, 3.8,
4.66, 1.387, 1.736,
4.056, 2.358, 2.07,
4.891, 1.393, 0.566,
3.662, 0.25, 1.744,
3.905, -0.749, 1.073,
2.585, 0.272, 2.505,
2.322, 0.419, 3.646,
1.744, 0.737, 1.804,
7.676, 2.1, 1.198,
7.457, 3.022, 0.385,
8.555, 1.167, 0.933,
9.232, 0.619, 1.734,
9.355, 1.03, -0.303,
8.921, 1.826, -1.066,
10.789, 1.367, -0.07,
11.352, 0.56, 0.612,
10.835, 2.302, 0.682,
11.708, 1.865, -1.158,
12.029, 3.005, -0.996,
13.04, 1.125, -1.019,
13.755, 1.775, -0.305,
13.695, 1.034, -2.022,
13.136, -0.003, -0.622,
11.168, 1.795, -2.571,
11.013, 0.691, -2.993,
10.457, 2.729, -2.8,
12.077, 2.106, -3.298,
9.322, -0.476, -0.629,
9.747, -1.293, 0.185,
8.695, -0.87, -1.734,
9.081, -0.26, -2.672,
8.54, -2.259, -2.038,
9.58, -2.666, -1.624,
7.12, -2.79, -1.68,
7.003, -3.882, -2.126,
6.773, -2.671, -0.222,
7.078, -3.7, 0.296,
7.258, -1.714, 0.295,
5.622, -2.596, 0.07,
6.149, -2.038, -2.393,
6.563, -0.948, -2.576,
8.789, -2.595, -3.498,
8.814, -1.84, -4.455,
9.039, -3.896, -3.649,
9.998, -4.257, -3.044,
9.213, -4.439, -5.004,
9.635, -3.601, -5.733,
10.362, -5.368, -5.148,
10.762, -5.554, -6.263,
11.388, -5.182, -4.551,
10.111, -6.488, -4.808,
7.831, -5.097, -5.245,
7.215, -5.663, -4.314,
7.344, -4.846, -6.46,
8.185, -5.251, -7.194,
6.039, -5.394, -6.815,
5.424, -5.934, -5.958,
5.029, -4.326, -7.188,
5.598, -3.545, -7.893,
4.874, -3.627, -6.236,
3.883, -4.767, -8.083,
3.509, -5.864, -7.803,
4.313, -4.917, -9.185,
2.67, -3.844, -8.025,
1.851, -4.238, -7.255,
2.922, -2.71, -7.769,
1.981, -3.77, -9.393,
1.818, -4.823, -9.939,
0.873, -3.359, -9.245,
2.784, -3.023, -10.42,
2.079, -3.106, -11.384,
2.831, -1.85, -10.218,
3.827, -3.479, -10.769,
6.246, -6.457, -7.903,
6.801, -6.201, -8.977,
5.859, -7.669, -7.551,
6.106, -8.022, -6.446,
5.918, -8.806, -8.452,
6.419, -8.545, -9.491,
6.677, -9.948, -7.747,
6.207, -10.409, -6.751,
6.552, -10.908, -8.455,
8.176, -9.565, -7.632,
8.538, -8.495, -7.254,
8.858, -10.451, -6.621,
8.196, -10.993, -5.784,
9.391, -11.431, -7.073,
9.816, -9.945, -6.106,
8.789, -9.713, -9.018,
8.866, -10.887, -9.265,
8.358, -9.316, -10.054,
9.947, -9.423, -8.895,
4.543, -9.275, -8.879,
3.654, -9.651, -8.1,
4.293, -9.259, -10.183,
4.438, -8.284, -10.848,
2.985, -9.682, -10.665,
2.786, -10.588, -9.916,
2.29, -8.809, -11.088,
3.02, -10.574, -11.897,
3.953, -10.662, -12.686,
1.885, -11.226, -12.06,
1.306, -11.693, -11.137,
1.649, -12.092, -13.195,
2.607, -12, -13.891,
1.739, -13.537, -12.685,
1.115, -14.042, -11.799,
2.846, -13.771, -12.291,
1.535, -14.515, -13.824,
2.565, -14.741, -14.74,
3.668, -14.926, -14.33,
2.385, -15.627, -15.79,
3.342, -15.961, -16.413,
1.173, -16.284, -15.914,
0.979, -17.172, -16.952,
1.921, -17.123, -17.665,
0.146, -16.067, -15.013,
-0.798, -16.772, -15.169,
0.326, -15.179, -13.969,
-0.06, -15.809, -13.036,
0.309, -11.751, -13.825,
-0.729, -11.638, -13.162,
0.274, -11.568, -15.129,
1.43, -11.664, -16.046,
1.942, -12.713, -16.279,
2.175, -10.752, -15.849,
0.853, -11.321, -17.404,
1.563, -10.614, -18.062,
0.815, -12.264, -18.144,
-0.519, -10.781, -17.224,
-1.117, -11.086, -18.216,
-0.445, -9.599, -17.385,
-0.963, -11.267, -15.83,
-1.637, -10.348, -15.503,
-1.888, -12.452, -16.009,
-1.626, -13.224, -16.917,
-2.921, -12.645, -15.243,
-2.964, -12.089, -14.2,
-3.94, -13.656, -15.383,
-3.422, -14.696, -15.658,
-5.011, -13.593, -14.262,
-5.787, -12.725, -14.505,
-6.055, -14.682, -14.48,
-7.033, -14.653, -15.172,
-5.696, -15.797, -14.749,
-6.631, -14.885, -13.445,
-4.372, -13.73, -12.898,
-5.212, -12.944, -12.551,
-4.428, -14.077, -11.749,
-3.254, -14.755, -12.847,
-2.961, -15.456, -11.916,
-2.205, -14.287, -13.162,
-3.578, -15.721, -13.482,
-4.73, -13.498, -16.707,
-5.057, -14.518, -17.309,
-5.081, -12.287, -17.099,
-4.615, -11.347, -16.557,
-5.773, -11.934, -18.31,
-5.59, -12.76, -19.153,
-7.264, -11.628, -18.19,
-7.917, -11.563, -19.188,
-8.022, -12.741, -17.476,
-9.194, -12.541, -17.663,
-7.933, -13.84, -17.946,
-8.04, -12.789, -16.285,
-7.454, -10.359, -17.505,
-6.764, -9.578, -18.022,
-5.075, -10.701, -18.909,
-3.984, -10.395, -18.43,
-5.646, -9.988, -19.871,
-6.245, -10.608, -20.693,
-4.974, -8.825, -20.438,
-3.797, -8.991, -20.54,
-5.409, -8.49, -21.878,
-4.727, -7.626, -22.349,
-6.533, -8.21, -22.173,
-5.135, -9.568, -22.906,
-3.977, -10.038, -23.044,
-6.134, -9.939, -23.582,
-5.281, -7.568, -19.603,
-4.615, -6.535, -19.751,
-6.316, -7.714, -18.797,
-7.149, -8.017, -19.594,
-6.836, -6.721, -17.911,
-6.54, -5.585, -18.091,
-8.371, -6.697, -18.139,
-8.989, -7.717, -18.067,
-8.956, -5.933, -17.433,
-8.823, -6.044, -19.426,
-8.07, -5.349, -20.17,
-10.03, -6.247, -19.71,
-6.582, -6.985, -16.415,
-6.58, -6.034, -15.624,
-6.418, -8.216, -15.973,
-5.421, -8.574, -16.509,
-6.242, -8.576, -14.61,
-6.487, -7.556, -14.06,
-7.266, -9.666, -14.234,
-6.731, -10.721, -14.116,
-8.089, -9.788, -15.093,
-8.189, -9.417, -13.06,
-9.335, -9.27, -13.363,
-8.397, -10.722, -12.278,
-9.311, -10.643, -11.497,
-8.901, -11.559, -12.981,
-7.618, -11.406, -11.679,
-7.662, -8.365, -12.092,
-8.581, -7.608, -12.049,
-7.867, -9.006, -11.106,
-6.522, -8.111, -11.879,
-4.884, -9.113, -14.196,
-4.399, -10.133, -14.719,
-4.259, -8.409, -13.23,
-4.094, -7.291, -13.598,
-3.001, -8.879, -12.673,
-2.645, -9.831, -13.282,
-1.869, -7.905, -12.626,
-0.865, -8.254, -12.079,
-2.11, -6.856, -12.114,
-1.187, -7.492, -13.878,
-1.039, -8.25, -14.83,
-0.754, -6.315, -13.941,
-3.187, -9.316, -11.197,
-4.06, -8.793, -10.485,
-2.371, -10.28, -10.827,
-1.533, -10.776, -11.494,
-2.329, -10.689, -9.402,
-2.949, -9.923, -8.748,
-2.698, -12.098, -8.984,
-2.693, -12.214, -7.794,
-4.112, -12.428, -9.442,
-4.614, -11.869, -10.367,
-4.792, -12.443, -8.453,
-4.358, -13.59, -9.601,
-1.72, -13.135, -9.543,
-0.714, -12.513, -9.348,
-1.255, -13.671, -10.513,
-2.048, -14.555, -9.173,
-2.384, -14.529, -8.018,
-1.052, -15.216, -9.013,
-2.821, -15.376, -9.58,
-0.882, -10.315, -8.987,
0.027, -10.386, -9.814,
-0.656, -9.837, -7.795,
-1.412, -9.943, -6.891,
0.68, -9.388, -7.419,
1.192, -10.451, -7.611,
0.943, -7.906, -7.859,
1.18, -6.922, -8.505,
1.536, -8.45, -8.744,
0.078, -6.922, -7.089,
0.464, -6.445, -5.834,
1.624, -6.537, -5.631,
-0.327, -5.564, -5.14,
0.065, -4.916, -4.235,
-1.555, -5.166, -5.663,
-2.339, -4.292, -4.936,
-1.781, -3.254, -4.943,
-1.983, -5.645, -6.911,
-2.723, -4.893, -7.442,
-1.171, -6.52, -7.603,
-1.264, -6.589, -8.784,
0.855, -9.5, -5.916,
-0.08, -9.754, -5.139,
2.122, -9.347, -5.575,
3.025, -9.821, -6.18,
2.571, -9.301, -4.203,
1.593, -8.918, -3.652,
3.256, -10.535, -3.567,
3.706, -10.577, -2.462,
2.292, -11.715, -3.559,
1.169, -11.824, -3.163,
2.266, -12.324, -4.593,
2.801, -12.547, -2.855,
4.411, -10.9, -4.343,
5.252, -10.099, -4.134,
3.567, -8.126, -4.186,
4.182, -7.848, -5.22,
3.653, -7.546, -3.016,
3.049, -7.752, -2.025,
4.627, -6.476, -2.785,
5.424, -6.719, -3.629,
3.948, -5.136, -2.485,
4.796, -4.363, -2.172,
3.381, -5.255, -1.445,
3.206, -4.579, -3.664,
4.084, -4.582, -4.461,
2.269, -5.301, -3.778,
2.656, -3.183, -3.55,
3.263, -2.173, -3.366,
2.421, -3.053, -4.712,
1.627, -2.996, -2.492,
0.714, -2.403, -2.961,
1.953, -2.53, -1.278,
3.244, -2.238, -1.005,
3.602, -1.127, -1.231,
3.492, -2.913, -0.059,
1.038, -2.378, -0.321,
0.682, -1.245, -0.389,
0.626, -3.157, 0.462,
5.46, -6.943, -1.587,
4.887, -7.504, -0.649,
6.76, -6.723, -1.644,
7.522, -6.422, -2.493,
7.59, -7.057, -0.501,
6.886, -6.748, 0.406,
8.16, -8.447, -0.502,
7.205, -9.168, -0.509,
8.702, -8.684, 0.538,
9.141, -8.856, -1.567,
10.099, -8.155, -1.696,
9.835, -10.143, -1.145,
9.175, -11.132, -0.988,
10.525, -10.086, -0.164,
10.653, -10.502, -1.951,
8.437, -9.067, -2.91,
7.49, -9.782, -2.76,
9.193, -9.783, -3.505,
8.267, -8.188, -3.694,
8.65, -5.98, -0.321,
9.225, -5.493, -1.289,
8.824, -5.59, 0.958,
9.062, -6.499, 1.687,
9.795, -4.553, 1.268,
10.874, -5.079, 1.309,
10.035, -3.739, 0.436,
9.74, -4.1, 2.708,
9.482, -4.847, 3.669,
10.024, -2.79, 2.873,
10.95, -2.364, 2.258,
10.072, -2.288, 4.249,
10.142, -3.158, 5.057,
11.191, -1.86, 4.346,
9.323, -1.003, 4.434,
9.043, -0.252, 3.504,
8.942, -0.779, 5.676,
9.986, -0.797, 6.246,
8.22, 0.359, 6.164,
8.462, 1.109, 5.279,
6.773, -0.074, 6.414,
6.035, -0.716, 5.744,
6.822, -0.735, 7.407,
5.895, 1.144, 6.725,
5.826, 2.119, 6.058,
5.914, 1.374, 7.891,
4.255, 0.52, 7.236,
3.322, 1.407, 5.921,
2.353, 0.804, 6.28,
3.904, 0.829, 5.072,
2.999, 2.468, 6.349,
8.727, 0.937, 7.503,
9.017, 0.307, 8.517,
8.82, 2.241, 7.459,
9.213, 2.743, 6.458,
9.172, 3.11, 8.539,
9.862, 2.569, 9.339,
10.09, 4.276, 8.091,
9.568, 5.124, 7.44,
10.422, 5.169, 9.28,
9.596, 5.514, 10.075,
10.745, 6.245, 8.848,
11.377, 4.925, 9.964,
11.38, 3.718, 7.512,
12.338, 3.663, 8.228,
11.522, 2.732, 6.847,
11.74, 4.568, 6.741,
7.84, 3.667, 9.077,
7.145, 4.427, 8.374,
7.492, 3.317, 10.297,
8.326, 3.394, 11.133,
6.275, 3.85, 10.863,
6.137, 4.886, 10.294,
5.317, 2.662, 10.98,
5.03, 2.215, 9.913,
4.211, 2.745, 11.424,
5.885, 1.567, 11.832,
6.567, 0.467, 11.424,
6.699, 0.056, 10.323,
6.889, -0.338, 12.484,
7.509, -1.303, 12.773,
6.43, 0.255, 13.631,
6.543, -0.167, 14.956,
6.789, -1.266, 15.335,
5.972, 0.652, 15.904,
5.916, 0.165, 16.987,
5.328, 1.848, 15.558,
4.91, 2.31, 16.563,
5.227, 2.281, 14.244,
4.111, 2.62, 14.026,
5.792, 1.467, 13.263,
6.383, 4.529, 12.225,
7.291, 4.469, 13.05,
5.26, 5.18, 12.547,
4.689, 5.754, 11.682,
5.053, 5.905, 13.758,
5.836, 5.513, 14.553,
5.375, 7.4, 13.523,
4.688, 7.897, 12.683,
6.48, 7.579, 13.097,
5.221, 8.199, 14.841,
4.121, 8.259, 15.292,
6.086, 7.907, 15.606,
5.513, 9.667, 14.566,
4.977, 10.074, 13.573,
6.654, 9.868, 14.26,
4.926, 10.562, 15.533,
4.364, 11.468, 14.996,
5.521, 11.021, 16.634,
6.753, 10.658, 16.913,
7.508, 11.049, 17.747,
7.529, 10.75, 16.009,
4.88, 11.836, 17.462,
5.561, 12.621, 18.049,
3.972, 12.565, 17.196,
3.618, 5.844, 14.257,
2.725, 6.298, 13.551,
3.418, 5.354, 15.474,
4.109, 4.679, 16.156,
2.081, 5.369, 16.083,
1.215, 5.521, 15.29,
1.671, 4.017, 16.571,
2.204, 3.611, 17.566,
0.566, 4.113, 17.02,
1.867, 3.082, 15.853,
2.088, 6.461, 17.172,
3.036, 6.657, 17.945,
1.06, 7.277, 17.176,
0.862, 7.739, 16.101,
0.839, 8.339, 18.139,
1.857, 8.52, 18.721,
0.682, 9.708, 17.537,
-0.022, 9.97, 16.608,
0.264, 10.505, 18.328,
1.988, 10.339, 17.143,
2.704, 10.88, 18.01,
2.346, 10.321, 15.947,
-0.412, 7.979, 18.957,
-1.492, 7.855, 18.387,
-0.256, 7.775, 20.262,
0.697, 8.398, 20.538,
-1.382, 7.479, 21.121,
-2.376, 7.463, 20.473,
-1.27, 6.23, 21.983,
-1.889, 5.926, 22.958,
-1.341, 4.959, 21.145,
-0.288, 4.384, 21.154,
-2.043, 4.156, 21.692,
-1.627, 5.054, 19.994,
-0.027, 6.225, 22.703,
0.363, 7.332, 22.753,
-1.693, 8.701, 22.013,
-1.083, 9.766, 21.958,
-2.741, 8.496, 22.791,
-3.433, 7.532, 22.757,
-3.289, 9.443, 23.727,
-2.285, 9.871, 24.191,
-4.218, 10.478, 23.115,
-4.779, 9.642, 22.469,
-4.449, 11.289, 22.26,
-4.425, 11.663, 24.041,
-3.436, 12.633, 24.16,
-3.072, 13.019, 23.096,
-3.59, 13.718, 25,
-2.981, 14.726, 24.854,
-4.752, 13.853, 25.74,
-4.882, 14.952, 26.565,
-4.505, 15.906, 25.975,
-5.753, 12.907, 25.638,
-6.842, 13.302, 25.909,
-5.582, 11.816, 24.794,
-6.621, 11.247, 24.701,
-4.023, 8.703, 24.859,
-4.612, 7.646, 24.676,
-3.893, 9.279, 26.038,
-3.252, 10.259, 26.209,
-4.46, 8.765, 27.282,
-5.422, 8.123, 26.989,
-3.442, 7.921, 28.05,
-3.387, 7.072, 27.197,
-2.265, 7.985, 28.231,
-4.023, 7.239, 29.139,
-3.48, 6.198, 29.311,
-4.896, 9.967, 28.116,
-4.334, 11.051, 27.91,
-5.879, 9.793, 28.985,
-6.628, 8.924, 28.681,
-6.338, 10.941, 29.801,
-6.193, 12.023, 29.32,
-7.804, 10.866, 30.155,
-8.398, 11.619, 29.438,
-8.165, 11.21, 31.242,
-8.458, 9.513, 29.963,
-9.227, 9.313, 29.015,
-8.155, 8.576, 30.861,
-8.256, 7.421, 30.587,
-8.654, 8.723, 31.934,
-5.432, 11.041, 31.034,
-5.059, 12.123, 31.482,
-5.063, 9.857, 31.521,
-5.412, 8.817, 31.074,
-4.167, 9.722, 32.653,
-4.579, 10.407, 33.54,
-4.013, 8.253, 33.113,
-3.51, 7.434, 32.411,
-3.147, 8.151, 34.37,
-3.674, 8.68, 35.311,
-2.055, 8.636, 34.469,
-2.997, 7.032, 34.778,
-5.348, 7.582, 33.349,
-5.657, 7.757, 34.497,
-5.286, 6.384, 33.268,
-6.425, 7.764, 32.86,
-2.766, 10.217, 32.234,
-2.316, 11.29, 32.61,
-2.138, 9.407, 31.409,
-2.817, 9.031, 30.515,
-0.822, 9.491, 30.87,
-0.12, 9.922, 31.737,
-0.435, 8.066, 30.359,
-0.517, 7.53, 29.295,
0.759, 8.179, 30.321,
-0.472, 7.039, 31.475,
0.383, 7.159, 32.569,
1.399, 7.767, 32.692,
0.37, 6.233, 33.596,
1.177, 6.238, 34.471,
-0.511, 5.178, 33.54,
-0.516, 4.266, 34.567,
0.459, 3.599, 34.47,
-1.374, 5.034, 32.473,
-1.954, 3.997, 32.477,
-1.353, 5.96, 31.441,
-1.265, 5.253, 30.486,
-0.505, 10.487, 29.782,
0.689, 10.763, 29.561,
-1.485, 11.062, 29.098,
-2.328, 11.603, 29.737,
-1.192, 12.036, 28.033,
-2.12, 12.737, 27.763,
-0.422, 12.797, 28.542,
-0.69, 11.349, 26.745,
-0.86, 10.138, 26.503,
-0.027, 12.148, 25.909,
0.58, 13.019, 26.449,
0.545, 11.716, 24.659,
-0.392, 11.243, 24.106,
1.014, 12.939, 23.83,
1.648, 12.576, 22.883,
1.842, 13.514, 24.476,
-0.062, 13.894, 23.394,
-0.705, 13.335, 22.557,
-0.661, 14.335, 24.325,
0.51, 15.037, 22.571,
1.424, 14.728, 21.864,
-0.294, 15.382, 21.75,
0.792, 16.279, 23.399,
0.706, 16.336, 24.592,
-0.008, 17.114, 23.089,
2.199, 16.761, 23.157,
2.925, 16.669, 24.107,
2.914, 16.388, 22.272,
2.127, 17.943, 22.968,
1.784, 10.801, 24.763,
2.707, 11.046, 25.541,
1.815, 9.763, 23.926,
1.092, 9.908, 23,
2.876, 8.863, 23.689,
3.787, 9.582, 23.971,
2.937, 7.557, 24.473,
2.523, 6.439, 24.358,
2.237, 7.87, 25.395,
4.404, 7.185, 24.738,
5.334, 7.997, 24.545,
4.631, 5.96, 25.185,
5.4, 5.871, 26.092,
4.399, 4.842, 24.847,
3.02, 8.55, 22.188,
2.117, 8.647, 21.378,
4.238, 8.205, 21.791,
5.223, 8.611, 22.319,
4.55, 7.858, 20.423,
3.58, 7.209, 20.189,
5.191, 8.961, 19.625,
4.589, 9.946, 19.932,
5.178, 8.858, 18.441,
6.603, 9.293, 19.951,
7.058, 10.602, 19.93,
6.577, 11.597, 20.373,
8.336, 10.618, 20.243,
9.177, 11.421, 20.493,
8.735, 9.368, 20.471,
7.671, 8.524, 20.293,
8.308, 7.521, 20.281,
5.431, 6.601, 20.43,
6.003, 6.203, 21.445,
5.506, 6.034, 19.243,
5.229, 6.59, 18.238,
6.318, 4.83, 19.048,
7.233, 4.925, 19.808,
5.559, 3.589, 19.402,
4.657, 3.157, 18.754,
5.041, 3.676, 20.478,
6.425, 2.402, 19.75,
7.664, 2.518, 19.86,
5.8, 1.317, 19.917,
6.854, 4.849, 17.626,
6.308, 5.49, 16.735,
7.988, 4.225, 17.434,
8.786, 3.886, 18.249,
8.63, 4.22, 16.109,
7.764, 4.336, 15.308,
9.623, 5.364, 16.092,
10.056, 5.717, 17.149,
10.802, 5.206, 15.157,
11.156, 6.186, 14.56,
11.178, 4.374, 14.383,
11.68, 5.082, 15.971,
8.858, 6.532, 15.727,
9.604, 7.373, 15.351,
9.098, 2.832, 15.784,
9.251, 1.917, 16.621,
9.242, 2.58, 14.475,
9.341, 3.42, 13.647,
9.632, 1.235, 14.063,
10.671, 1.173, 14.66,
9.085, 0.243, 14.434,
10.022, 1.196, 12.612,
9.845, 2.077, 11.78,
10.653, 0.086, 12.297,
11.173, -0.565, 13.149,
11.084, -0.272, 10.958,
10.513, 0.422, 10.187,
12.535, -0.126, 10.663,
13.159, -0.865, 11.364,
12.788, -0.406, 9.164,
13.382, 0.482, 8.614,
12.21, -0.915, 8.25,
13.662, -1.225, 9.288,
13.031, 1.298, 10.955,
12.858, 1.71, 12.066,
12.954, 2.26, 10.249,
14.225, 1.153, 10.984,
10.558, -1.703, 10.813,
10.641, -2.535, 11.714,
9.848, -1.95, 9.693,
10.275, -1.705, 8.617,
9.291, -3.336, 9.653,
10.372, -3.765, 9.929,
7.98, -3.157, 10.438,
8.256, -3.018, 11.59,
7.15, -2.413, 10.018,
7.258, -4.317, 10.666,
7.074, -4.85, 9.632,
9.164, -3.853, 8.263,
8.948, -3.135, 7.278,
9.31, -5.157, 8.073,
9.579, -6.182, 9.109,
9.672, -5.511, 10.092,
9.548, -7.079, 9.912,
10.165, -7.283, 8.259,
11.307, -6.938, 8.111,
10.401, -8.426, 8.535,
9.409, -7.245, 6.97,
10.108, -7.717, 6.119,
8.472, -7.982, 6.976,
9.097, -5.759, 6.762,
10.036, -5.405, 6.121,
7.61, -5.581, 6.409,
6.738, -5.704, 7.295,
7.308, -5.313, 5.121,
7.828, -6.21, 4.54,
5.91, -5.235, 4.722,
5.305, -5.372, 5.732,
5.39, -3.936, 4.056,
5.12, -4.107, 2.905,
4.091, -3.547, 4.687,
3.634, -3.857, 5.737,
3.3, -3.852, 3.846,
4.069, -2.351, 4.733,
6.418, -2.896, 3.87,
7.207, -2.984, 4.76,
5.949, -1.802, 3.821,
6.986, -2.974, 2.824,
5.625, -6.235, 3.572,
6.423, -6.442, 2.658,
4.442, -6.782, 3.604,
4.053, -6.841, 4.71,
3.985, -7.71, 2.594,
4.706, -7.63, 1.655,
4.018, -9.144, 3.133,
3.266, -9.254, 4.047,
3.796, -10.026, 2.359,
5.38, -9.58, 3.636,
6.43, -9.747, 2.757,
6.246, -10.514, 1.866,
7.682, -10.135, 3.213,
8.636, -10.511, 2.612,
7.888, -10.366, 4.55,
8.895, -10.896, 4.898,
6.842, -10.185, 5.439,
7.077, -10.784, 6.435,
5.619, -9.785, 4.993,
4.907, -9.685, 5.934,
2.583, -7.379, 2.135,
1.738, -6.947, 2.917,
2.31, -7.627, 0.847,
2.829, -8.623, 0.46,
0.943, -7.418, 0.356,
0.35, -8.012, 1.198,
0.67, -6.029, -0.165,
1.539, -5.94, -0.971,
0.916, -5.28, 0.723,
-0.33, -5.947, -0.803,
0.628, -8.431, -0.75,
1.522, -8.885, -1.467,
-0.65, -8.729, -0.829,
-1.566, -8.878, -0.09,
-1.099, -9.604, -1.961,
-0.351, -10.035, -2.775,
-1.585, -10.633, -1.584,
-2.34, -8.872, -2.516,
-3.158, -8.313, -1.772,
-2.48, -8.807, -3.826,
-2.2, -9.811, -4.399,
-3.656, -8.06, -4.326,
-3.263, -6.942, -4.252,
-4.545, -8.702, -3.848,
-3.948, -8.379, -5.775,
-3.327, -9.212, -6.439,
-4.966, -7.688, -6.265,
-5.971, -7.375, -5.723,
-5.375, -7.813, -7.676,
-4.345, -8.127, -8.173,
-6.666, -8.618, -7.779,
-7.288, -8.785, -6.773,
-7.695, -8.034, -8.697,
-8.349, -7.192, -8.139,
-7.411, -7.353, -9.63,
-8.611, -8.802, -8.805,
-6.328, -10.047, -8.261,
-5.176, -10.308, -8.133,
-6.785, -10.735, -7.385,
-6.914, -10.543, -9.176,
-5.436, -6.397, -8.219,
-5.845, -5.462, -7.493,
-4.996, -6.219, -9.435,
-4.715, -6.991, -10.28,
-5.018, -4.924, -10.104,
-5.587, -4.192, -9.367,
-3.623, -4.411, -10.417,
-3.094, -5.146, -9.637,
-2.688, -4.564, -11.157,
-3.663, -2.941, -10.788,
-4.387, -2.145, -10.281,
-3.784, -2.994, -11.974,
-2.383, -2.187, -10.559,
-1.509, -2.215, -11.432,
-2.251, -1.529, -9.504,
-5.83, -5.067, -11.414,
-5.514, -5.952, -12.213,
-6.886, -4.28, -11.598,
-6.415, -3.197, -11.615,
-7.708, -4.405, -12.812,
-7.531, -5.37, -13.479,
-9.114, -4.826, -12.438,
-9.737, -3.995, -11.844,
-9.294, -5.679, -11.622,
-10.105, -5.007, -13.55,
-10.646, -3.893, -14.173,
-10.209, -2.798, -14.181,
-11.556, -4.003, -15.205,
-12.332, -3.281, -15.74,
-11.964, -5.252, -15.628,
-12.886, -5.317, -16.661,
-12.296, -5.59, -17.648,
-11.449, -6.375, -15.026,
-11.947, -7.402, -15.365,
-10.523, -6.256, -14,
-9.965, -7.292, -14.103,
-7.633, -3.152, -13.66,
-8.013, -2.057, -13.244,
-7.126, -3.281, -14.884,
-6.15, -3.957, -14.893,
-6.997, -2.134, -15.788,
-6.339, -1.346, -15.189,
-5.994, -2.318, -16.896,
-5.527, -1.272, -17.242,
-5.085, -2.974, -16.493,
-6.458, -2.707, -17.928,
-8.35, -1.86, -16.453,
-8.725, -2.643, -17.299,
-8.998, -0.805, -16.008,
-8.38, -0.199, -15.212,
-10.283, -0.411, -16.542,
-11.01, -1.328, -16.765,
-10.873, 0.811, -15.815,
-10.617, 1.953, -16.024,
-12.32, 1.01, -16.31,
-12.552, 1.963, -17.006,
-13.153, 1.235, -15.475,
-12.877, 0.158, -16.949,
-10.854, 0.691, -14.308,
-11.442, 1.625, -13.839,
-9.854, 0.726, -13.665,
-11.626, -0.523, -13.774,
-12.11, -1.345, -14.495,
-11.538, -1.142, -12.756,
-12.678, -0.033, -13.446,
-10.031, 0.019, -18.012,
-10.672, -0.447, -18.936,
-9.094, 0.937, -18.147,
-8.662, 1.597, -17.267,
-8.629, 1.504, -19.366,
-8.976, 0.778, -20.248,
-9.018, 2.978, -19.57,
-9.251, 3.326, -20.692,
-10.407, 3.285, -19.092,
-10.557, 3.677, -17.974,
-11.191, 2.439, -19.415,
-10.856, 4.217, -19.709,
-8.048, 3.779, -18.875,
-8.368, 4.905, -19.044,
-7.105, 1.426, -19.271,
-6.589, 0.98, -18.261,
-6.398, 1.841, -20.281,
-6.863, 2.366, -21.593,
-7.847, 1.953, -22.137,
-6.877, 3.49, -22.003,
-5.806, 1.715, -22.483,
-6.292, 0.656, -22.773,
-5.451, 2.025, -23.589,
-4.53, 1.911, -21.708,
-3.63, 1.199, -22.032,
-4.061, 2.98, -21.976,
-4.94, 1.742, -20.255,
-4.63, 0.638, -19.937,
-4.331, 2.721, -19.284,
-3.188, 2.474, -18.854,
-5.023, 3.781, -18.87,
-5.55, 4.223, -19.834,
-4.422, 4.684, -17.892,
-3.267, 4.431, -17.834,
-4.499, 6.151, -18.305,
-4.593, 6.944, -17.419,
-3.478, 6.456, -18.848,
-5.753, 6.453, -19.121,
-5.712, 7.651, -19.221,
-6.889, 6.401, -18.764,
-5.384, 6.404, -20.616,
-4.229, 6.801, -20.879,
-6.228, 5.976, -21.418,
-5.024, 4.573, -16.493,
-4.49, 5.181, -15.547,
-6.135, 3.848, -16.32,
-6.434, 2.925, -16.993,
-6.683, 3.827, -14.979,
-5.756, 4.144, -14.312,
-7.751, 4.842, -14.637,
-7.314, 5.586, -13.81,
-8.117, 6.082, -15.448,
-8.591, 5.88, -16.528,
-7.378, 7.009, -15.624,
-9, 6.715, -14.932,
-9.071, 4.106, -14.312,
-9.138, 3.405, -15.268,
-10.092, 4.71, -14.492,
-9.143, 4.082, -12.796,
-8.197, 4.579, -12.267,
-9.489, 2.988, -12.475,
-10.095, 4.728, -12.443,
-6.891, 2.397, -14.518,
-7.525, 1.529, -15.129,
-6.305, 2.137, -13.311,
-5.22, 2.472, -12.976,
-6.45, 0.765, -12.8,
-7.361, 0.203, -13.3,
-5.064, 0.073, -12.86,
-4.565, 0.343, -13.911,
-4.364, 0.378, -11.941,
-5.18, -1.112, -12.842,
-6.981, 0.762, -11.379,
-6.727, 1.685, -10.62,
-7.714, -0.264, -10.976,
-7.443, -1.319, -11.424,
-8.168, -0.319, -9.578,
-8.086, 0.687, -8.964,
-9.677, -0.598, -9.494,
-10.164, -1.109, -8.531,
-10.538, 0.59, -9.867,
-10.391, 1.44, -10.69,
-11.641, 0.177, -10.108,
-10.811, 1.175, -8.858,
-9.939, -1.702, -10.402,
-9.96, -1.265, -11.493,
-7.398, -1.487, -8.929,
-7.012, -2.401, -9.662,
-7.177, -1.432, -7.615,
-6.695, -0.395, -7.312,
-6.543, -2.471, -6.882,
-7.171, -3.289, -7.487,
-5.104, -2.362, -6.569,
-4.833, -2.352, -7.729,
-4.656, -3.332, -6.04,
-4.388, -1.24, -5.899,
-4.309, -1.513, -4.738,
-4.835, -0.136, -5.848,
-3.13, -1.005, -6.788,
-2.799, -1.978, -7.395,
-3.253, -0.045, -7.485,
-1.934, -1.006, -6.074,
-2.113, -0.57, -4.98,
-0.68, -0.887, -6.402,
-0.28, -0.779, -7.664,
-0.152, -1.56, -8.545,
0.082, 0.263, -8.099,
0.221, -0.883, -5.393,
0.153, -0.214, -4.413,
0.821, -1.892, -5.531,
-7.351, -2.851, -5.619,
-8.018, -2.072, -4.989,
-7.284, -4.138, -5.327,
-6.335, -4.749, -5.672,
-7.9, -4.75, -4.143,
-8.313, -3.862, -3.477,
-9.056, -5.603, -4.481,
-9.796, -4.924, -5.136,
-8.811, -6.485, -5.249,
-10.036, -6.18, -3.474,
-11.126, -6.205, -3.97,
-9.688, -7.629, -3.141,
-10.653, -8.251, -3.497,
-9.596, -7.98, -1.998,
-8.818, -8.254, -3.68,
-10.146, -5.352, -2.191,
-10.114, -4.167, -2.121,
-11.236, -5.671, -1.8,
-9.449, -5.715, -1.289,
-6.673, -5.433, -3.515,
-5.961, -6.216, -4.122,
-6.297, -5.017, -2.331,
-6.45, -3.879, -2.051,
-5.071, -5.491, -1.717,
-5.144, -6.622, -2.074,
-3.989, -4.41, -2.003,
-3.863, -4.195, -3.166,
-4.252, -3.352, -1.514,
-2.651, -4.675, -1.356,
-2.252, -5.661, -1.888,
-2.688, -4.679, -0.166,
-1.671, -3.524, -1.522,
-1.072, -3.454, -2.597,
-1.476, -2.698, -0.611,
-5.23, -5.689, -0.219,
-5.967, -4.974, 0.466,
-4.484, -6.651, 0.256,
-4.734, -7.669, -0.306,
-4.378, -6.994, 1.66,
-5.025, -6.296, 2.359,
-4.842, -8.437, 1.919,
-5.901, -8.987, 1.811,
-4.209, -9.246, 1.303,
-4.58, -8.818, 3.363,
-5.372, -8.2, 4.35,
-6.194, -7.35, 4.375,
-5.184, -8.477, 5.679,
-6.177, -8.634, 6.319,
-4.188, -9.384, 6.03,
-4.035, -9.635, 7.377,
-3.268, -10.528, 7.508,
-3.379, -10.003, 5.093,
-2.992, -11.109, 5.297,
-3.579, -9.698, 3.744,
-3.315, -10.652, 3.084,
-2.879, -6.828, 2.026,
-1.977, -7.466, 1.464,
-2.593, -5.919, 2.934,
-3.19, -4.9, 2.845,
-1.204, -5.661, 3.358,
-0.497, -6.256, 2.62,
-0.956, -4.162, 3.247,
-1.245, -3.753, 2.163,
-1.594, -3.553, 4.048,
0.419, -3.645, 3.504,
0.668, -3.79, 4.661,
1.29, -4.024, 2.789,
0.48, -2.126, 3.367,
0.48, -1.557, 2.251,
0.531, -1.499, 4.536,
-0.266, -1.362, 5.411,
1.544, -1.275, 5.116,
-0.973, -6.11, 4.794,
-1.782, -5.867, 5.719,
0.165, -6.725, 5.053,
1.079, -6.115, 4.619,
0.447, -7.093, 6.446,
0.069, -6.13, 7.04,
0.013, -8.493, 6.841,
-0.324, -9.43, 7.524,
-0.9, -7.992, 7.436,
0.822, -9.605, 6.247,
1.822, -10.304, 6.861,
2.054, -10.497, 8.009,
2.34, -11.243, 5.995,
2.914, -12.228, 6.331,
1.688, -11.162, 4.799,
1.858, -11.887, 3.616,
2.533, -12.863, 3.546,
1.043, -11.555, 2.541,
1.117, -12.327, 1.64,
0.074, -10.536, 2.619,
-0.722, -10.822, 1.786,
-0.088, -9.821, 3.798,
-0.961, -9.027, 3.849,
0.718, -10.131, 4.915,
1.919, -6.86, 6.717,
2.759, -6.752, 5.845,
2.201, -6.731, 8.001,
1.35, -6.712, 8.827,
3.59, -6.597, 8.48,
4.333, -6.93, 7.616,
3.916, -5.27, 9.142,
5.084, -5.081, 9.098,
3.275, -4.081, 8.435,
2.312, -3.614, 8.978,
2.74, -4.317, 7.401,
3.988, -3.119, 8.475,
3.438, -5.379, 10.482,
4.191, -4.79, 11.181,
3.734, -7.732, 9.505,
2.763, -7.973, 10.236,
4.859, -8.438, 9.487,
5.701, -8.439, 8.654,
4.934, -9.514, 10.53,
3.88, -9.905, 10.93,
5.442, -10.799, 9.991,
4.715, -11.326, 9.202,
5.619, -11.668, 10.797,
6.827, -10.786, 9.402,
7.216, -11.728, 8.704,
7.592, -9.736, 9.664,
8.106, -8.942, 10.382,
8.614, -10.268, 9.336,
5.69, -8.888, 11.698,
6.596, -8.061, 11.455,
5.268, -9.144, 12.935,
4.499, -10.001, 13.234,
5.935, -8.517, 14.089,
6.923, -8.578, 13.439,
5.294, -7.171, 14.433,
5.495, -6.723, 15.522,
4.124, -7.278, 14.249,
5.788, -5.973, 13.652,
5.119, -4.932, 13.546,
6.98, -6.061, 13.06,
7.483, -6.166, 11.994,
7.769, -5.498, 13.756,
5.982, -9.441, 15.298,
5.007, -9.703, 16,
7.967, -8.857, 14.94,
8.649, -8.19, 14.233,
9.093, -9.317, 15.831,
8.618, -10.039, 16.649,
10.187, -10.099, 15.036,
10.631, -9.61, 14.042,
11.438, -10.384, 15.884,
12.436, -10.775, 15.344,
11.263, -11.145, 16.794,
11.951, -9.448, 16.43,
9.705, -11.497, 14.578,
9.2, -12.185, 15.417,
8.869, -11.396, 13.729,
10.826, -12.386, 14.022,
10.464, -12.649, 12.909,
12.001, -12.263, 13.84,
10.747, -13.464, 14.54,
9.672, -8.074, 16.653,
9.533, -7.966, 17.849,
10.384, -7.074, 16.113,
11.14, -7.137, 15.197,
10.748, -5.788, 16.892,
10.145, -4.99, 17.555,
10.507, -5.155, 15.9,
11.744, -5.896, 18.096,
11.726, -6.832, 18.901,
12.603, -4.867, 18.184,
12.698, -4.083, 17.294,
13.605, -4.736, 19.262,
13.884, -5.803, 19.716,
14.924, -4.212, 18.693,
15.486, -3.772, 19.657,
15.155, -3.283, 17.969,
15.553, -5.171, 17.677,
14.927, -6.246, 17.331,
16.706, -4.903, 17.163,
13.051, -3.783, 20.319,
12.368, -2.793, 19.996,
13.315, -4.079, 21.588,
14.188, -4.814, 21.924,
12.84, -3.175, 22.635,
13.629, -2.289, 22.489,
11.331, -2.954, 22.522,
10.827, -3.555, 21.618,
10.412, -3.048, 23.284,
11.219, -1.795, 22.22,
13.01, -3.61, 24.106,
13.813, -4.561, 24.375,
12.171, -2.737, 24.733,
12.639, -1.662, 24.508,
11.749, -2.477, 26.151,
11.412, -1.324, 26.112,
11.19, -3.612, 27.043,
10.314, -2.998, 26.431,
10.867, -2.902, 28.015,
10.414, -4.752, 26.511,
10.836, -5.68, 25.525,
11.265, -5.443, 24.438,
9.781, -6.473, 25.301,
9.19, -6.047, 24.349,
8.803, -6.099, 26.11,
9.216, -5.082, 26.909,
8.094, -5.266, 27.363,
12.601, -2.602, 27.275,
13.24, -1.483, 27.569,
11.943, -3.843, 27.298,
13.092, -4.183, 27.469,
11.663, -5.225, 27.936,
12.309, -5.692, 28.828,
10.118, -5.195, 28.1,
9.969, -6.189, 28.77,
9.65, -4.393, 29.305,
9.096, -3.346, 29.529,
8.758, -5.023, 29.822,
10.439, -4.361, 30.212,
9.563, -4.524, 26.94,
8.779, -3.632, 27.246,
11.832, -6.35, 26.764,
12.709, -6.247, 25.909,
10.956, -7.43, 26.668,
10.531, -7.994, 27.625,
11.042, -8.483, 25.541,
12.074, -8.34, 24.961,
11.198, -9.918, 26.091,
10.235, -10.262, 26.708,
11.383, -10.976, 24.989,
10.562, -11.83, 25.187,
12.419, -11.581, 24.944,
11.269, -10.868, 23.802,
12.416, -10.074, 27.008,
13.461, -9.816, 26.481,
12.489, -9.523, 28.069,
12.604, -11.501, 27.529,
11.728, -11.724, 28.321,
12.679, -12.568, 26.985,
13.625, -11.509, 28.163,
9.771, -8.445, 24.627,
8.646, -8.264, 25.107,
9.993, -8.635, 23.316,
11.117, -8.813, 22.957,
8.936, -8.52, 22.254,
9.523, -7.463, 22.164,
9.503, -9.276, 21.495,
7.959, -9.747, 22.173,
8.383, -10.895, 22.446,
6.667, -9.372, 21.768,
6.11, -8.724, 22.603,
5.44, -10.292, 21.53,
5.703, -11.361, 21.066,
4.768, -10.663, 22.826,
3.732, -11.253, 22.755,
5.686, -11.444, 23.769,
6.414, -12.298, 23.343,
4.898, -12.133, 24.359,
6.31, -11.015, 24.699,
4.35, -9.492, 23.51,
5.013, -9.337, 24.479,
4.467, -9.714, 20.419,
4.89, -9.247, 19.358,
3.055, -9.646, 20.399,
2.198, -9.843, 21.198,
2.709, -9.092, 19.073,
2.793, -7.923, 19.302,
3.746, -9.998, 18.278,
3.424, -10.159, 17.141,
3.642, -11.151, 18.606,
5.296, -9.46, 18.478,
5.963, -10.429, 18.227,
5.415, -8.642, 17.61,
5.848, -8.828, 19.871,
5.522, -8.14, 20.818,
5.618, -7.685, 19.465,
7.196, -8.104, 19.663,
7.45, -7.7, 18.574,
8.138, -7.658, 20.593,
7.997, -7.819, 21.917,
7.579, -7.697, 23.052,
7.473, -6.726, 21.809,
9.297, -7.016, 20.258,
8.891, -6.201, 19.482,
10.165, -6.348, 20.734,
1.118, -8.749, 18.482,
0.094, -9.074, 19.173,
1.164, -8.628, 17.114,
0.486, -9.347, 16.616,
-0.447, -9.933, 16.118,
1.133, -9.697, 15.656,
0.678, -9.696, 17.972,
-0.174, -10.555, 18.134,
1.418, -10.65, 18.003,
-0.169, -8.442, 18.162,
-0.546, -7.553, 18.9,
-1.328, -8.777, 18.016,
0.3, -7.8, 16.896,
-0.67, -7.73, 16.184,
0.376, -6.455, 16.71,
0.064, -5.967, 17.915,
1.083, -6.37, 15.011,
2.011, -7.099, 14.973,
0.427, -5.645, 13.913,
-0.224, -4.869, 14.533,
1.523, -4.974, 13.067,
2.673, -4.884, 12.76,
1.691, -4.126, 13.903,
1.075, -4.677, 11.649,
1.024, -5.595, 10.791,
0.781, -3.504, 11.345,
-0.404, -6.566, 13.028,
0.105, -7.611, 12.591,
-1.629, -6.204, 12.668,
-1.757, -5.031, 12.575,
-2.469, -7.056, 11.812,
-1.963, -8.128, 11.663,
-3.8, -7.285, 12.521,
-4.424, -6.284, 12.464,
-3.534, -7.86, 13.534,
-4.671, -8.39, 11.981,
-4.233, -9.525, 11.765,
-5.954, -8.078, 11.751,
-6.336, -8.741, 10.834,
-6.954, -7.619, 12.196,
-2.657, -6.505, 10.405,
-2.077, -5.482, 10.046,
-3.428, -7.163, 9.534,
-3.745, -8.305, 9.606,
-3.552, -6.715, 8.189,
-2.432, -6.39, 7.968,
-4.13, -7.471, 7.483,
-4.437, -5.531, 7.907,
-5.383, -5.212, 8.609,
-4.14, -4.886, 6.784,
-3.018, -4.554, 6.599,
-4.93, -3.799, 6.267,
-5.88, -3.697, 6.972,
-4.139, -2.512, 6.162,
-3.753, -2.127, 7.222,
-3.176, -2.51, 5.463,
-4.954, -1.322, 5.718,
-5.444, -1.438, 4.643,
-5.682, -0.799, 6.497,
-4.019, 0.198, 5.56,
-3.153, -0.018, 4.039,
-2.222, 0.379, 4.668,
-3.015, -1.055, 3.479,
-3.937, 0.788, 3.654,
-5.479, -4.209, 4.88,
-4.739, -4.646, 3.983,
-6.781, -4.07, 4.726,
-7.556, -3.632, 5.497,
-7.446, -4.316, 3.454,
-6.747, -4.95, 2.744,
-8.86, -4.889, 3.586,
-9.234, -4.857, 4.719,
-9.618, -4.342, 2.848,
-8.96, -6.389, 3.339,
-8.597, -7.06, 4.258,
-10.442, -6.785, 3.233,
-10.511, -7.973, 3.426,
-11.1, -6.739, 2.231,
-11.168, -6.496, 4.138,
-8.208, -6.803, 2.074,
-8.823, -7.802, 1.806,
-7.138, -7.29, 1.943,
-8.566, -6.121, 1.157,
-7.648, -2.977, 2.741,
-8.049, -1.998, 3.379,
-7.403, -2.94, 1.443,
-6.345, -3.214, 0.993,
-7.654, -1.651, 0.78,
-8.738, -1.423, 1.22,
-6.443, -0.762, 1.018,
-6.625, 0.357, 0.661,
-5.996, -0.786, 2.122,
-5.373, -1.234, 0.254,
-4.389, -1.055, 0.879,
-8.099, -1.72, -0.655,
-7.908, -2.709, -1.369,
-8.762, -0.651, -1.09,
-9.249, 0.167, -0.386,
-9.243, -0.484, -2.448,
-9.077, -1.454, -3.103,
-10.713, -0.011, -2.415,
-10.958, 1.008, -1.841,
-10.976, 0.313, -3.539,
-11.743, -1.016, -1.937,
-11.597, -1.334, -0.799,
-13.098, -0.319, -1.954,
-13.278, 0.792, -1.539,
-13.865, -0.946, -1.277,
-13.676, -0.225, -3.003,
-11.728, -2.261, -2.82,
-11.999, -3.121, -2.034,
-11.079, -2.422, -3.811,
-12.78, -2.329, -3.402,
-8.469, 0.733, -2.976,
-8.486, 1.713, -2.239,
-7.94, 0.736, -4.169,
-8.448, 0.04, -4.983,
-7.157, 1.879, -4.66,
-6.044, 1.47, -4.574,
-7.592, 2.847, -4.123,
-7.486, 2.043, -6.158,
-8.073, 1.18, -6.803,
-7.122, 3.206, -6.656,
-7.12, 4.162, -5.952,
-7.201, 3.677, -7.986,
-7.453, 2.715, -8.625,
-8.218, 4.811, -8.145,
-8.057, 5.869, -7.611,
-8.373, 5.147, -9.624,
-7.649, 6.051, -9.932,
-9.404, 5.727, -9.837,
-8.571, 4.061, -10.067,
-9.586, 4.343, -7.657,
-10.17, 3.351, -7.976,
-10.445, 5.155, -7.88,
-9.703, 4.334, -6.462,
-5.81, 4.231, -8.355,
-5.11, 4.845, -7.539,
-5.373, 3.966, -9.576,
-6.048, 3.665, -10.497,
-4.122, 4.53, -10.017,
-4.282, 5.596, -9.508,
-2.869, 3.741, -9.734,
-1.825, 4.302, -9.83,
-3.017, 3.22, -8.674,
-2.65, 2.63, -10.488,
-2.064, 2.948, -11.463,
-4.195, 4.968, -11.488,
-4.859, 4.419, -12.356,
-3.426, 6.009, -11.695,
-3.421, 6.905, -10.914,
-3.252, 6.614, -12.992,
-4.265, 6.401, -13.576,
-3.451, 8.121, -12.837,
-2.758, 8.81, -12.146,
-4.511, 8.449, -12.383,
-3.374, 8.817, -14.175,
-4.448, 8.753, -15.052,
-5.569, 8.776, -14.653,
-4.4, 9.386, -16.278,
-5.367, 9.87, -16.777,
-3.259, 10.08, -16.622,
-3.199, 10.722, -17.851,
-2.061, 10.82, -18.157,
-2.171, 10.146, -15.774,
-1.58, 11.172, -15.862,
-2.217, 9.514, -14.545,
-1.342, 9.812, -13.803,
-1.872, 6.283, -13.555,
-0.838, 6.413, -12.911,
-1.866, 5.821, -14.809,
-2.576, 6.43, -15.535,
-0.6, 5.493, -15.464,
0.299, 5.351, -14.703,
-0.672, 4.125, -16.168,
-1.347, 4.196, -17.146,
0.378, 3.965, -16.723,
-0.876, 2.966, -15.2,
0.149, 2.552, -14.763,
-1.565, 3.334, -14.298,
-1.659, 1.869, -15.813,
-1.012, 1.662, -16.795,
-2.802, 2.148, -16.011,
-1.839, 0.731, -14.909,
-1.823, 0.886, -13.731,
-2.046, -0.488, -15.407,
-2.081, -0.624, -16.727,
-2.547, 0.194, -17.457,
-2.038, -1.439, -17.59,
-2.208, -1.538, -14.629,
-2.64, -1.427, -13.53,
-2.014, -2.707, -14.69,
-0.232, 6.56, -16.478,
-1.064, 6.83, -17.359,
0.931, 7.156, -16.314,
1.817, 6.734, -15.66,
1.463, 8.133, -17.269,
0.666, 8.831, -17.816,
2.501, 9.017, -16.548,
2.639, 9.9, -17.35,
3.645, 8.733, -16.344,
2.03, 9.688, -15.317,
1.402, 10.924, -15.362,
1.564, 11.748, -16.205,
0.948, 11.553, -14.208,
0.633, 12.701, -14.229,
1.117, 10.944, -12.981,
1.103, 11.768, -12.123,
1.737, 9.698, -12.91,
2.551, 9.824, -12.052,
2.183, 9.086, -14.071,
3.271, 8.669, -13.852,
2.207, 7.33, -18.337,
3.453, 7.331, -18.274,
1.616, 6.557, -19.217,
0.671, 7.054, -19.744,
2.355, 5.742, -20.172,
2.775, 4.726, -19.721,
1.538, 5.456, -20.996,
3.434, 6.468, -20.955,
4.41, 7.074, -20.476;
	charges = 
-0.4157,
0.2719,
-0.0237,
0.088,
0.0342,
0.0241,
0.0241,
0.0018,
0.044,
0.044,
-0.2737,
-0.0536,
0.0684,
0.0684,
0.0684,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.3479,
0.2747,
-0.24,
0.1426,
-0.0094,
0.0362,
0.0362,
0.0187,
0.0103,
0.0103,
-0.0479,
0.0621,
0.0621,
-0.0143,
0.1135,
0.1135,
-0.3854,
0.34,
0.34,
0.34,
0.7341,
-0.5894,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0275,
0.1123,
-0.005,
0.0339,
0.0339,
-0.1415,
-0.1638,
0.2062,
-0.3418,
0.3412,
0.138,
-0.2601,
0.1572,
-0.1134,
0.1417,
-0.1972,
0.1447,
-0.2387,
0.17,
0.1243,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.24,
0.1426,
-0.0094,
0.0362,
0.0362,
0.0187,
0.0103,
0.0103,
-0.0479,
0.0621,
0.0621,
-0.0143,
0.1135,
0.1135,
-0.3854,
0.34,
0.34,
0.34,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0275,
0.1123,
-0.005,
0.0339,
0.0339,
-0.1415,
-0.1638,
0.2062,
-0.3418,
0.3412,
0.138,
-0.2601,
0.1572,
-0.1134,
0.1417,
-0.1972,
0.1447,
-0.2387,
0.17,
0.1243,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0249,
0.0843,
0.2117,
0.0352,
0.0352,
-0.6546,
0.4275,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0031,
0.085,
-0.0036,
0.0171,
0.0171,
-0.0645,
0.0352,
0.0352,
0.6951,
-0.6086,
-0.9407,
0.4251,
0.4251,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0188,
0.0881,
-0.0462,
0.0402,
0.0402,
-0.0266,
-0.3811,
0.3649,
0.2057,
0.1392,
-0.5727,
0.1292,
0.1147,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0597,
0.0869,
0.1303,
0.0187,
-0.3204,
0.0882,
0.0882,
0.0882,
-0.043,
0.0236,
0.0236,
-0.066,
0.0186,
0.0186,
0.0186,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0188,
0.0881,
-0.0462,
0.0402,
0.0402,
-0.0266,
-0.3811,
0.3649,
0.2057,
0.1392,
-0.5727,
0.1292,
0.1147,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0397,
0.1105,
0.056,
-0.0173,
-0.0173,
0.0136,
-0.0425,
-0.0425,
0.8054,
-0.8188,
-0.8188,
0.5366,
-0.5819,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.24,
0.1426,
-0.0094,
0.0362,
0.0362,
0.0187,
0.0103,
0.0103,
-0.0479,
0.0621,
0.0621,
-0.0143,
0.1135,
0.1135,
-0.3854,
0.34,
0.34,
0.34,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0024,
0.0978,
-0.0343,
0.0295,
0.0295,
0.0118,
-0.1256,
0.133,
-0.1704,
0.143,
-0.1072,
0.1297,
-0.1704,
0.143,
-0.1256,
0.133,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0031,
0.085,
-0.0036,
0.0171,
0.0171,
-0.0645,
0.0352,
0.0352,
0.6951,
-0.6086,
-0.9407,
0.4251,
0.4251,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0024,
0.0978,
-0.0343,
0.0295,
0.0295,
0.0118,
-0.1256,
0.133,
-0.1704,
0.143,
-0.1072,
0.1297,
-0.1704,
0.143,
-0.1256,
0.133,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0397,
0.1105,
0.056,
-0.0173,
-0.0173,
0.0136,
-0.0425,
-0.0425,
0.8054,
-0.8188,
-0.8188,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0237,
0.088,
0.0342,
0.0241,
0.0241,
0.0018,
0.044,
0.044,
-0.2737,
-0.0536,
0.0684,
0.0684,
0.0684,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0275,
0.1123,
-0.005,
0.0339,
0.0339,
-0.1415,
-0.1638,
0.2062,
-0.3418,
0.3412,
0.138,
-0.2601,
0.1572,
-0.1134,
0.1417,
-0.1972,
0.1447,
-0.2387,
0.17,
0.1243,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.2637,
0.156,
-0.0007,
0.0327,
0.0327,
0.039,
0.0285,
0.0285,
0.0486,
0.0687,
0.0687,
-0.5295,
0.3456,
0.8076,
-0.8627,
0.4478,
0.4478,
-0.8627,
0.4478,
0.4478,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0237,
0.088,
0.0342,
0.0241,
0.0241,
0.0018,
0.044,
0.044,
-0.2737,
-0.0536,
0.0684,
0.0684,
0.0684,
0.5973,
-0.5679,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.24,
0.1426,
-0.0094,
0.0362,
0.0362,
0.0187,
0.0103,
0.0103,
-0.0479,
0.0621,
0.0621,
-0.0143,
0.1135,
0.1135,
-0.3854,
0.34,
0.34,
0.34,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0249,
0.0843,
0.2117,
0.0352,
0.0352,
-0.6546,
0.4275,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0397,
0.1105,
0.056,
-0.0173,
-0.0173,
0.0136,
-0.0425,
-0.0425,
0.8054,
-0.8188,
-0.8188,
0.5366,
-0.5819,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.24,
0.1426,
-0.0094,
0.0362,
0.0362,
0.0187,
0.0103,
0.0103,
-0.0479,
0.0621,
0.0621,
-0.0143,
0.1135,
0.1135,
-0.3854,
0.34,
0.34,
0.34,
0.7341,
-0.5894,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0031,
0.085,
-0.0036,
0.0171,
0.0171,
-0.0645,
0.0352,
0.0352,
0.6951,
-0.6086,
-0.9407,
0.4251,
0.4251,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0031,
0.085,
-0.0036,
0.0171,
0.0171,
-0.0645,
0.0352,
0.0352,
0.6951,
-0.6086,
-0.9407,
0.4251,
0.4251,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.24,
0.1426,
-0.0094,
0.0362,
0.0362,
0.0187,
0.0103,
0.0103,
-0.0479,
0.0621,
0.0621,
-0.0143,
0.1135,
0.1135,
-0.3854,
0.34,
0.34,
0.34,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.4157,
0.2719,
-0.0597,
0.0869,
0.1303,
0.0187,
-0.3204,
0.0882,
0.0882,
0.0882,
-0.043,
0.0236,
0.0236,
-0.066,
0.0186,
0.0186,
0.0186,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0597,
0.0869,
0.1303,
0.0187,
-0.3204,
0.0882,
0.0882,
0.0882,
-0.043,
0.0236,
0.0236,
-0.066,
0.0186,
0.0186,
0.0186,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.2637,
0.156,
-0.0007,
0.0327,
0.0327,
0.039,
0.0285,
0.0285,
0.0486,
0.0687,
0.0687,
-0.5295,
0.3456,
0.8076,
-0.8627,
0.4478,
0.4478,
-0.8627,
0.4478,
0.4478,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0237,
0.088,
0.0342,
0.0241,
0.0241,
0.0018,
0.044,
0.044,
-0.2737,
-0.0536,
0.0684,
0.0684,
0.0684,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0275,
0.1123,
-0.005,
0.0339,
0.0339,
-0.1415,
-0.1638,
0.2062,
-0.3418,
0.3412,
0.138,
-0.2601,
0.1572,
-0.1134,
0.1417,
-0.1972,
0.1447,
-0.2387,
0.17,
0.1243,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.2637,
0.156,
-0.0007,
0.0327,
0.0327,
0.039,
0.0285,
0.0285,
0.0486,
0.0687,
0.0687,
-0.5295,
0.3456,
0.8076,
-0.8627,
0.4478,
0.4478,
-0.8627,
0.4478,
0.4478,
0.7341,
-0.5894,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0249,
0.0843,
0.2117,
0.0352,
0.0352,
-0.6546,
0.4275,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.24,
0.1426,
-0.0094,
0.0362,
0.0362,
0.0187,
0.0103,
0.0103,
-0.0479,
0.0621,
0.0621,
-0.0143,
0.1135,
0.1135,
-0.3854,
0.34,
0.34,
0.34,
0.7341,
-0.5894,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0188,
0.0881,
-0.0462,
0.0402,
0.0402,
-0.0266,
-0.3811,
0.3649,
0.2057,
0.1392,
-0.5727,
0.1292,
0.1147,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0249,
0.0843,
0.2117,
0.0352,
0.0352,
-0.6546,
0.4275,
0.5973,
-0.5679,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0024,
0.0978,
-0.0343,
0.0295,
0.0295,
0.0118,
-0.1256,
0.133,
-0.1704,
0.143,
-0.1072,
0.1297,
-0.1704,
0.143,
-0.1256,
0.133,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0397,
0.1105,
0.056,
-0.0173,
-0.0173,
0.0136,
-0.0425,
-0.0425,
0.8054,
-0.8188,
-0.8188,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0597,
0.0869,
0.1303,
0.0187,
-0.3204,
0.0882,
0.0882,
0.0882,
-0.043,
0.0236,
0.0236,
-0.066,
0.0186,
0.0186,
0.0186,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.5163,
0.2936,
0.0397,
0.1105,
0.056,
-0.0173,
-0.0173,
0.0136,
-0.0425,
-0.0425,
0.8054,
-0.8188,
-0.8188,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0597,
0.0869,
0.1303,
0.0187,
-0.3204,
0.0882,
0.0882,
0.0882,
-0.043,
0.0236,
0.0236,
-0.066,
0.0186,
0.0186,
0.0186,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.2637,
0.156,
-0.0007,
0.0327,
0.0327,
0.039,
0.0285,
0.0285,
0.0486,
0.0687,
0.0687,
-0.5295,
0.3456,
0.8076,
-0.8627,
0.4478,
0.4478,
-0.8627,
0.4478,
0.4478,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0397,
0.1105,
0.056,
-0.0173,
-0.0173,
0.0136,
-0.0425,
-0.0425,
0.8054,
-0.8188,
-0.8188,
0.5366,
-0.5819,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0031,
0.085,
-0.0036,
0.0171,
0.0171,
-0.0645,
0.0352,
0.0352,
0.6951,
-0.6086,
-0.9407,
0.4251,
0.4251,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0275,
0.1123,
-0.005,
0.0339,
0.0339,
-0.1415,
-0.1638,
0.2062,
-0.3418,
0.3412,
0.138,
-0.2601,
0.1572,
-0.1134,
0.1417,
-0.1972,
0.1447,
-0.2387,
0.17,
0.1243,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0597,
0.0869,
0.1303,
0.0187,
-0.3204,
0.0882,
0.0882,
0.0882,
-0.043,
0.0236,
0.0236,
-0.066,
0.0186,
0.0186,
0.0186,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
0.0337,
0.0823,
-0.1825,
0.0603,
0.0603,
0.0603,
0.5973,
-0.5679,
-0.4157,
0.2719,
0.0188,
0.0881,
-0.0462,
0.0402,
0.0402,
-0.0266,
-0.3811,
0.3649,
0.2057,
0.1392,
-0.5727,
0.1292,
0.1147,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0597,
0.0869,
0.1303,
0.0187,
-0.3204,
0.0882,
0.0882,
0.0882,
-0.043,
0.0236,
0.0236,
-0.066,
0.0186,
0.0186,
0.0186,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0389,
0.1007,
0.3654,
0.0043,
-0.2438,
0.0642,
0.0642,
0.0642,
-0.6761,
0.4102,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.2637,
0.156,
-0.0007,
0.0327,
0.0327,
0.039,
0.0285,
0.0285,
0.0486,
0.0687,
0.0687,
-0.5295,
0.3456,
0.8076,
-0.8627,
0.4478,
0.4478,
-0.8627,
0.4478,
0.4478,
0.7341,
-0.5894,
-0.2548,
0.0192,
0.0391,
0.0391,
0.0189,
0.0213,
0.0213,
-0.007,
0.0253,
0.0253,
-0.0266,
0.0641,
0.5896,
-0.5748,
-0.5163,
0.2936,
0.0381,
0.088,
-0.0303,
-0.0122,
-0.0122,
0.7994,
-0.8014,
-0.8014,
0.5366,
-0.5819,
-0.4157,
0.2719,
0.0143,
0.1048,
-0.2041,
0.0797,
0.0797,
0.713,
-0.5931,
-0.9191,
0.4196,
0.4196,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0237,
0.088,
0.0342,
0.0241,
0.0241,
0.0018,
0.044,
0.044,
-0.2737,
-0.0536,
0.0684,
0.0684,
0.0684,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0249,
0.0843,
0.2117,
0.0352,
0.0352,
-0.6546,
0.4275,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0518,
0.0922,
-0.1102,
0.0457,
0.0457,
0.3531,
-0.0361,
-0.4121,
0.1,
0.1,
0.1,
-0.4121,
0.1,
0.1,
0.1,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0875,
0.0969,
0.2985,
-0.0297,
-0.3192,
0.0791,
0.0791,
0.0791,
-0.3192,
0.0791,
0.0791,
0.0791,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0249,
0.0843,
0.2117,
0.0352,
0.0352,
-0.6546,
0.4275,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0014,
0.0876,
-0.0152,
0.0295,
0.0295,
-0.0011,
-0.1906,
0.1699,
-0.2341,
0.1656,
0.3226,
-0.5579,
0.3992,
-0.2341,
0.1656,
-0.1906,
0.1699,
0.5973,
-0.5679,
-0.3479,
0.2747,
-0.2637,
0.156,
-0.0007,
0.0327,
0.0327,
0.039,
0.0285,
0.0285,
0.0486,
0.0687,
0.0687,
-0.5295,
0.3456,
0.8076,
-0.8627,
0.4478,
0.4478,
-0.8627,
0.4478,
0.4478,
0.7341,
-0.5894,
-0.4157,
0.2719,
-0.0024,
0.0978,
-0.0343,
0.0295,
0.0295,
0.0118,
-0.1256,
0.133,
-0.1704,
0.143,
-0.1072,
0.1297,
-0.1704,
0.143,
-0.1256,
0.133,
0.5973,
-0.5679,
-0.4157,
0.2719,
-0.0252,
0.0698,
0.0698,
0.5973,
-0.5679;
	radii = 
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
2,
1.908,
1.387,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.1,
1.1,
1.824,
0.6,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.409,
1.824,
0.6,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.1,
1.1,
1.824,
0.6,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.409,
1.824,
0.6,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.387,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.824,
0.6,
1.908,
1.359,
1.824,
1.908,
1.409,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.824,
0.6,
1.908,
1.359,
1.824,
1.908,
1.409,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.1,
1.1,
1.824,
0.6,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
2,
1.908,
1.387,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.409,
1.824,
0.6,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
1.824,
0.6,
1.908,
1.824,
0.6,
0.6,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
2,
1.908,
1.387,
1.387,
1.387,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.1,
1.1,
1.824,
0.6,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.387,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.1,
1.1,
1.824,
0.6,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.1,
1.1,
1.824,
0.6,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
1.824,
0.6,
1.908,
1.824,
0.6,
0.6,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
2,
1.908,
1.387,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.409,
1.824,
0.6,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
1.824,
0.6,
1.908,
1.824,
0.6,
0.6,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.387,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.1,
1.1,
1.824,
0.6,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.824,
0.6,
1.908,
1.359,
1.824,
1.908,
1.409,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.387,
1.721,
0,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
1.824,
0.6,
1.908,
1.824,
0.6,
0.6,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.409,
1.824,
0.6,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.824,
0.6,
1.908,
1.359,
1.824,
1.908,
1.409,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.908,
1.487,
1.487,
1.487,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
1.824,
0.6,
1.908,
1.824,
0.6,
0.6,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
1.908,
1.387,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.6612,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
2,
1.908,
1.387,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.387,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.487,
1.487,
1.487,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.387,
1.387,
1.721,
0,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.721,
0,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.487,
1.487,
1.908,
1.387,
1.387,
1.824,
0.6,
1.908,
1.824,
0.6,
0.6,
1.824,
0.6,
0.6,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.908,
1.487,
1.487,
1.908,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.459,
1.908,
1.6612,
1.824,
0.6,
1.908,
1.387,
1.387,
1.908,
1.6612;
	epsilon = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	mass = 
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
32.06,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
14.01,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
14.01,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
14.01,
1.008,
12.01,
1.008,
14.01,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
14.01,
1.008,
12.01,
1.008,
14.01,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
32.06,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
14.01,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
12.01,
14.01,
1.008,
1.008,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
32.06,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
12.01,
14.01,
1.008,
1.008,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
32.06,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
14.01,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
12.01,
14.01,
1.008,
1.008,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
14.01,
1.008,
12.01,
1.008,
14.01,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
12.01,
14.01,
1.008,
1.008,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
14.01,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
14.01,
1.008,
12.01,
1.008,
14.01,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
12.01,
14.01,
1.008,
1.008,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
16,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
32.06,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
1.008,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
16,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
12.01,
1.008,
1.008,
14.01,
1.008,
12.01,
14.01,
1.008,
1.008,
14.01,
1.008,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
12.01,
1.008,
1.008,
12.01,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
1.008,
12.01,
16,
14.01,
1.008,
12.01,
1.008,
1.008,
12.01,
16;
	surfaceaccessibility = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
	hydrophobicityscale = 
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.108,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
0.112,
0.0362,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
0.112,
0.0362,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.112,
0.0362,
-0.0134,
-0.0397,
0.112,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.112,
0.0362,
-0.0134,
-0.0397,
0.112,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.108,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
0.112,
0.0362,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
-0.0134,
0.112,
0.0362,
0.0362,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.108,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
-0.0134,
0.112,
0.0362,
0.0362,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.108,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
0.112,
0.0362,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
-0.0134,
0.112,
0.0362,
0.0362,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.112,
0.0362,
-0.0134,
-0.0397,
0.112,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
-0.0134,
0.112,
0.0362,
0.0362,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
0.112,
0.0362,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.112,
0.0362,
-0.0134,
-0.0397,
0.112,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
-0.0134,
0.112,
0.0362,
0.0362,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.0403,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.108,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.0403,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.0362,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.105,
-0.0397,
-0.0397,
0.112,
0.0362,
-0.0134,
0.112,
0.0362,
0.0362,
0.112,
0.0362,
0.0362,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.105,
-0.0397,
-0.0397,
-0.0134,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
-0.0397,
-0.0134,
0.0403,
0.112,
0.0362,
-0.105,
-0.0397,
-0.0397,
-0.0134,
0.0403;
	particlenames = 
"MN",
"MH",
"MCA",
"MHA",
"MCB",
"MHB2",
"MHB3",
"MCG",
"MHG2",
"MHG3",
"MSD",
"MCE",
"MHE1",
"MHE2",
"MHE3",
"MC",
"MO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"KN",
"KH",
"KCA",
"KHA",
"KCB",
"KHB2",
"KHB3",
"KCG",
"KHG2",
"KHG3",
"KCD",
"KHD2",
"KHD3",
"KCE",
"KHE2",
"KHE3",
"KNZ",
"KHZ1",
"KHZ2",
"KHZ3",
"KC",
"KO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"WN",
"WH",
"WCA",
"WHA",
"WCB",
"WHB2",
"WHB3",
"WCG",
"WCD1",
"WHD1",
"WNE1",
"WHE1",
"WCE2",
"WCZ2",
"WHZ2",
"WCH2",
"WHH2",
"WCZ3",
"WHZ3",
"WCE3",
"WHE3",
"WCD2",
"WC",
"WO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"KN",
"KH",
"KCA",
"KHA",
"KCB",
"KHB2",
"KHB3",
"KCG",
"KHG2",
"KHG3",
"KCD",
"KHD2",
"KHD3",
"KCE",
"KHE2",
"KHE3",
"KNZ",
"KHZ1",
"KHZ2",
"KHZ3",
"KC",
"KO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"WN",
"WH",
"WCA",
"WHA",
"WCB",
"WHB2",
"WHB3",
"WCG",
"WCD1",
"WHD1",
"WNE1",
"WHE1",
"WCE2",
"WCZ2",
"WHZ2",
"WCH2",
"WHH2",
"WCZ3",
"WHZ3",
"WCE3",
"WHE3",
"WCD2",
"WC",
"WO",
"SN",
"SH",
"SCA",
"SHA",
"SCB",
"SHB2",
"SHB3",
"SOG",
"SHG",
"SC",
"SO",
"QN",
"QH",
"QCA",
"QHA",
"QCB",
"QHB2",
"QHB3",
"QCG",
"QHG2",
"QHG3",
"QCD",
"QOE1",
"QNE2",
"QHE21",
"QHE22",
"QC",
"QO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"HN",
"HH",
"HCA",
"HHA",
"HCB",
"HHB2",
"HHB3",
"HCG",
"HND1",
"HHD1",
"HCE1",
"HHE1",
"HNE2",
"HCD2",
"HHD2",
"HC",
"HO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"IN",
"IH",
"ICA",
"IHA",
"ICB",
"IHB",
"ICG2",
"IHG21",
"IHG22",
"IHG23",
"ICG1",
"IHG12",
"IHG13",
"ICD1",
"IHD11",
"IHD12",
"IHD13",
"IC",
"IO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"HN",
"HH",
"HCA",
"HHA",
"HCB",
"HHB2",
"HHB3",
"HCG",
"HND1",
"HHD1",
"HCE1",
"HHE1",
"HNE2",
"HCD2",
"HHD2",
"HC",
"HO",
"EN",
"EH",
"ECA",
"EHA",
"ECB",
"EHB2",
"EHB3",
"ECG",
"EHG2",
"EHG3",
"ECD",
"EOE1",
"EOE2",
"EC",
"EO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"KN",
"KH",
"KCA",
"KHA",
"KCB",
"KHB2",
"KHB3",
"KCG",
"KHG2",
"KHG3",
"KCD",
"KHD2",
"KHD3",
"KCE",
"KHE2",
"KHE3",
"KNZ",
"KHZ1",
"KHZ2",
"KHZ3",
"KC",
"KO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"FN",
"FH",
"FCA",
"FHA",
"FCB",
"FHB2",
"FHB3",
"FCG",
"FCD1",
"FHD1",
"FCE1",
"FHE1",
"FCZ",
"FHZ",
"FCE2",
"FHE2",
"FCD2",
"FHD2",
"FC",
"FO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"QN",
"QH",
"QCA",
"QHA",
"QCB",
"QHB2",
"QHB3",
"QCG",
"QHG2",
"QHG3",
"QCD",
"QOE1",
"QNE2",
"QHE21",
"QHE22",
"QC",
"QO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"FN",
"FH",
"FCA",
"FHA",
"FCB",
"FHB2",
"FHB3",
"FCG",
"FCD1",
"FHD1",
"FCE1",
"FHE1",
"FCZ",
"FHZ",
"FCE2",
"FHE2",
"FCD2",
"FHD2",
"FC",
"FO",
"EN",
"EH",
"ECA",
"EHA",
"ECB",
"EHB2",
"EHB3",
"ECG",
"EHG2",
"EHG3",
"ECD",
"EOE1",
"EOE2",
"EC",
"EO",
"MN",
"MH",
"MCA",
"MHA",
"MCB",
"MHB2",
"MHB3",
"MCG",
"MHG2",
"MHG3",
"MSD",
"MCE",
"MHE1",
"MHE2",
"MHE3",
"MC",
"MO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"WN",
"WH",
"WCA",
"WHA",
"WCB",
"WHB2",
"WHB3",
"WCG",
"WCD1",
"WHD1",
"WNE1",
"WHE1",
"WCE2",
"WCZ2",
"WHZ2",
"WCH2",
"WHH2",
"WCZ3",
"WHZ3",
"WCE3",
"WHE3",
"WCD2",
"WC",
"WO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"RN",
"RH",
"RCA",
"RHA",
"RCB",
"RHB2",
"RHB3",
"RCG",
"RHG2",
"RHG3",
"RCD",
"RHD2",
"RHD3",
"RNE",
"RHE",
"RCZ",
"RNH1",
"RHH11",
"RHH12",
"RNH2",
"RHH21",
"RHH22",
"RC",
"RO",
"MN",
"MH",
"MCA",
"MHA",
"MCB",
"MHB2",
"MHB3",
"MCG",
"MHG2",
"MHG3",
"MSD",
"MCE",
"MHE1",
"MHE2",
"MHE3",
"MC",
"MO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"KN",
"KH",
"KCA",
"KHA",
"KCB",
"KHB2",
"KHB3",
"KCG",
"KHG2",
"KHG3",
"KCD",
"KHD2",
"KHD3",
"KCE",
"KHE2",
"KHE3",
"KNZ",
"KHZ1",
"KHZ2",
"KHZ3",
"KC",
"KO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"SN",
"SH",
"SCA",
"SHA",
"SCB",
"SHB2",
"SHB3",
"SOG",
"SHG",
"SC",
"SO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"EN",
"EH",
"ECA",
"EHA",
"ECB",
"EHB2",
"EHB3",
"ECG",
"EHG2",
"EHG3",
"ECD",
"EOE1",
"EOE2",
"EC",
"EO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"KN",
"KH",
"KCA",
"KHA",
"KCB",
"KHB2",
"KHB3",
"KCG",
"KHG2",
"KHG3",
"KCD",
"KHD2",
"KHD3",
"KCE",
"KHE2",
"KHE3",
"KNZ",
"KHZ1",
"KHZ2",
"KHZ3",
"KC",
"KO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"QN",
"QH",
"QCA",
"QHA",
"QCB",
"QHB2",
"QHB3",
"QCG",
"QHG2",
"QHG3",
"QCD",
"QOE1",
"QNE2",
"QHE21",
"QHE22",
"QC",
"QO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"QN",
"QH",
"QCA",
"QHA",
"QCB",
"QHB2",
"QHB3",
"QCG",
"QHG2",
"QHG3",
"QCD",
"QOE1",
"QNE2",
"QHE21",
"QHE22",
"QC",
"QO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"KN",
"KH",
"KCA",
"KHA",
"KCB",
"KHB2",
"KHB3",
"KCG",
"KHG2",
"KHG3",
"KCD",
"KHD2",
"KHD3",
"KCE",
"KHE2",
"KHE3",
"KNZ",
"KHZ1",
"KHZ2",
"KHZ3",
"KC",
"KO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"IN",
"IH",
"ICA",
"IHA",
"ICB",
"IHB",
"ICG2",
"IHG21",
"IHG22",
"IHG23",
"ICG1",
"IHG12",
"IHG13",
"ICD1",
"IHD11",
"IHD12",
"IHD13",
"IC",
"IO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"IN",
"IH",
"ICA",
"IHA",
"ICB",
"IHB",
"ICG2",
"IHG21",
"IHG22",
"IHG23",
"ICG1",
"IHG12",
"IHG13",
"ICD1",
"IHD11",
"IHD12",
"IHD13",
"IC",
"IO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"RN",
"RH",
"RCA",
"RHA",
"RCB",
"RHB2",
"RHB3",
"RCG",
"RHG2",
"RHG3",
"RCD",
"RHD2",
"RHD3",
"RNE",
"RHE",
"RCZ",
"RNH1",
"RHH11",
"RHH12",
"RNH2",
"RHH21",
"RHH22",
"RC",
"RO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"MN",
"MH",
"MCA",
"MHA",
"MCB",
"MHB2",
"MHB3",
"MCG",
"MHG2",
"MHG3",
"MSD",
"MCE",
"MHE1",
"MHE2",
"MHE3",
"MC",
"MO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"WN",
"WH",
"WCA",
"WHA",
"WCB",
"WHB2",
"WHB3",
"WCG",
"WCD1",
"WHD1",
"WNE1",
"WHE1",
"WCE2",
"WCZ2",
"WHZ2",
"WCH2",
"WHH2",
"WCZ3",
"WHZ3",
"WCE3",
"WHE3",
"WCD2",
"WC",
"WO",
"RN",
"RH",
"RCA",
"RHA",
"RCB",
"RHB2",
"RHB3",
"RCG",
"RHG2",
"RHG3",
"RCD",
"RHD2",
"RHD3",
"RNE",
"RHE",
"RCZ",
"RNH1",
"RHH11",
"RHH12",
"RNH2",
"RHH21",
"RHH22",
"RC",
"RO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"SN",
"SH",
"SCA",
"SHA",
"SCB",
"SHB2",
"SHB3",
"SOG",
"SHG",
"SC",
"SO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"KN",
"KH",
"KCA",
"KHA",
"KCB",
"KHB2",
"KHB3",
"KCG",
"KHG2",
"KHG3",
"KCD",
"KHD2",
"KHD3",
"KCE",
"KHE2",
"KHE3",
"KNZ",
"KHZ1",
"KHZ2",
"KHZ3",
"KC",
"KO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"HN",
"HH",
"HCA",
"HHA",
"HCB",
"HHB2",
"HHB3",
"HCG",
"HND1",
"HHD1",
"HCE1",
"HHE1",
"HNE2",
"HCD2",
"HHD2",
"HC",
"HO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"SN",
"SH",
"SCA",
"SHA",
"SCB",
"SHB2",
"SHB3",
"SOG",
"SHG",
"SC",
"SO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"FN",
"FH",
"FCA",
"FHA",
"FCB",
"FHB2",
"FHB3",
"FCG",
"FCD1",
"FHD1",
"FCE1",
"FHE1",
"FCZ",
"FHZ",
"FCE2",
"FHE2",
"FCD2",
"FHD2",
"FC",
"FO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"EN",
"EH",
"ECA",
"EHA",
"ECB",
"EHB2",
"EHB3",
"ECG",
"EHG2",
"EHG3",
"ECD",
"EOE1",
"EOE2",
"EC",
"EO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"IN",
"IH",
"ICA",
"IHA",
"ICB",
"IHB",
"ICG2",
"IHG21",
"IHG22",
"IHG23",
"ICG1",
"IHG12",
"IHG13",
"ICD1",
"IHD11",
"IHD12",
"IHD13",
"IC",
"IO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"EN",
"EH",
"ECA",
"EHA",
"ECB",
"EHB2",
"EHB3",
"ECG",
"EHG2",
"EHG3",
"ECD",
"EOE1",
"EOE2",
"EC",
"EO",
"IN",
"IH",
"ICA",
"IHA",
"ICB",
"IHB",
"ICG2",
"IHG21",
"IHG22",
"IHG23",
"ICG1",
"IHG12",
"IHG13",
"ICD1",
"IHD11",
"IHD12",
"IHD13",
"IC",
"IO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"RN",
"RH",
"RCA",
"RHA",
"RCB",
"RHB2",
"RHB3",
"RCG",
"RHG2",
"RHG3",
"RCD",
"RHD2",
"RHD3",
"RNE",
"RHE",
"RCZ",
"RNH1",
"RHH11",
"RHH12",
"RNH2",
"RHH21",
"RHH22",
"RC",
"RO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"EN",
"EH",
"ECA",
"EHA",
"ECB",
"EHB2",
"EHB3",
"ECG",
"EHG2",
"EHG3",
"ECD",
"EOE1",
"EOE2",
"EC",
"EO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"QN",
"QH",
"QCA",
"QHA",
"QCB",
"QHB2",
"QHB3",
"QCG",
"QHG2",
"QHG3",
"QCD",
"QOE1",
"QNE2",
"QHE21",
"QHE22",
"QC",
"QO",
"WN",
"WH",
"WCA",
"WHA",
"WCB",
"WHB2",
"WHB3",
"WCG",
"WCD1",
"WHD1",
"WNE1",
"WHE1",
"WCE2",
"WCZ2",
"WHZ2",
"WCH2",
"WHH2",
"WCZ3",
"WHZ3",
"WCE3",
"WHE3",
"WCD2",
"WC",
"WO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"IN",
"IH",
"ICA",
"IHA",
"ICB",
"IHB",
"ICG2",
"IHG21",
"IHG22",
"IHG23",
"ICG1",
"IHG12",
"IHG13",
"ICD1",
"IHD11",
"IHD12",
"IHD13",
"IC",
"IO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"AN",
"AH",
"ACA",
"AHA",
"ACB",
"AHB1",
"AHB2",
"AHB3",
"AC",
"AO",
"HN",
"HH",
"HCA",
"HHA",
"HCB",
"HHB2",
"HHB3",
"HCG",
"HND1",
"HHD1",
"HCE1",
"HHE1",
"HNE2",
"HCD2",
"HHD2",
"HC",
"HO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"IN",
"IH",
"ICA",
"IHA",
"ICB",
"IHB",
"ICG2",
"IHG21",
"IHG22",
"IHG23",
"ICG1",
"IHG12",
"IHG13",
"ICD1",
"IHD11",
"IHD12",
"IHD13",
"IC",
"IO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"TN",
"TH",
"TCA",
"THA",
"TCB",
"THB",
"TCG2",
"THG21",
"THG22",
"THG23",
"TOG1",
"THG1",
"TC",
"TO",
"RN",
"RH",
"RCA",
"RHA",
"RCB",
"RHB2",
"RHB3",
"RCG",
"RHG2",
"RHG3",
"RCD",
"RHD2",
"RHD3",
"RNE",
"RHE",
"RCZ",
"RNH1",
"RHH11",
"RHH12",
"RNH2",
"RHH21",
"RHH22",
"RC",
"RO",
"PN",
"PCD",
"PHD2",
"PHD3",
"PCG",
"PHG2",
"PHG3",
"PCB",
"PHB2",
"PHB3",
"PCA",
"PHA",
"PC",
"PO",
"DN",
"DH",
"DCA",
"DHA",
"DCB",
"DHB2",
"DHB3",
"DCG",
"DOD1",
"DOD2",
"DC",
"DO",
"NN",
"NH",
"NCA",
"NHA",
"NCB",
"NHB2",
"NHB3",
"NCG",
"NOD1",
"NND2",
"NHD21",
"NHD22",
"NC",
"NO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"MN",
"MH",
"MCA",
"MHA",
"MCB",
"MHB2",
"MHB3",
"MCG",
"MHG2",
"MHG3",
"MSD",
"MCE",
"MHE1",
"MHE2",
"MHE3",
"MC",
"MO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"SN",
"SH",
"SCA",
"SHA",
"SCB",
"SHB2",
"SHB3",
"SOG",
"SHG",
"SC",
"SO",
"LN",
"LH",
"LCA",
"LHA",
"LCB",
"LHB2",
"LHB3",
"LCG",
"LHG",
"LCD1",
"LHD11",
"LHD12",
"LHD13",
"LCD2",
"LHD21",
"LHD22",
"LHD23",
"LC",
"LO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO",
"VN",
"VH",
"VCA",
"VHA",
"VCB",
"VHB",
"VCG1",
"VHG11",
"VHG12",
"VHG13",
"VCG2",
"VHG21",
"VHG22",
"VHG23",
"VC",
"VO",
"SN",
"SH",
"SCA",
"SHA",
"SCB",
"SHB2",
"SHB3",
"SOG",
"SHG",
"SC",
"SO",
"YN",
"YH",
"YCA",
"YHA",
"YCB",
"YHB2",
"YHB3",
"YCG",
"YCD1",
"YHD1",
"YCE1",
"YHE1",
"YCZ",
"YOH",
"YHH",
"YCE2",
"YHE2",
"YCD2",
"YHD2",
"YC",
"YO",
"RN",
"RH",
"RCA",
"RHA",
"RCB",
"RHB2",
"RHB3",
"RCG",
"RHG2",
"RHG3",
"RCD",
"RHD2",
"RHD3",
"RNE",
"RHE",
"RCZ",
"RNH1",
"RHH11",
"RHH12",
"RNH2",
"RHH21",
"RHH22",
"RC",
"RO",
"FN",
"FH",
"FCA",
"FHA",
"FCB",
"FHB2",
"FHB3",
"FCG",
"FCD1",
"FHD1",
"FCE1",
"FHE1",
"FCZ",
"FHZ",
"FCE2",
"FHE2",
"FCD2",
"FHD2",
"FC",
"FO",
"GN",
"GH",
"GCA",
"GHA2",
"GHA3",
"GC",
"GO";
	resnames = 
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"LYS",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"GLU",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"GLN",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"TRP",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"ALA",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"HIS",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"ILE",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"THR",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"PRO",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASP",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"ASN",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"MET",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"LEU",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"VAL",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"SER",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"TYR",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"ARG",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"PHE",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY",
"GLY";
	resids = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
2,
2,
2,
2,
2,
2,
2,
2,
2,
2,
2,
2,
2,
2,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
3,
4,
4,
4,
4,
4,
4,
4,
4,
4,
4,
4,
4,
5,
5,
5,
5,
5,
5,
5,
5,
5,
5,
5,
5,
5,
5,
6,
6,
6,
6,
6,
6,
6,
6,
6,
6,
6,
6,
6,
6,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
7,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
8,
9,
9,
9,
9,
9,
9,
9,
9,
9,
9,
9,
9,
9,
9,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
12,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
13,
14,
14,
14,
14,
14,
14,
14,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
15,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
20,
20,
20,
20,
20,
20,
20,
20,
20,
20,
20,
20,
21,
21,
21,
21,
21,
21,
21,
21,
21,
21,
21,
21,
21,
21,
22,
22,
22,
22,
22,
22,
22,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
23,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
24,
25,
25,
25,
25,
25,
25,
25,
25,
25,
25,
25,
25,
25,
25,
26,
26,
26,
26,
26,
26,
26,
26,
26,
26,
26,
26,
26,
26,
27,
27,
27,
27,
27,
27,
27,
27,
27,
27,
27,
27,
27,
27,
28,
28,
28,
28,
28,
28,
28,
29,
29,
29,
29,
29,
29,
29,
29,
29,
29,
29,
29,
29,
29,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
30,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
31,
32,
32,
32,
32,
32,
32,
32,
32,
32,
32,
32,
32,
32,
32,
32,
33,
33,
33,
33,
33,
33,
33,
33,
33,
33,
33,
33,
33,
33,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
34,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
35,
36,
36,
36,
36,
36,
36,
36,
37,
37,
37,
37,
37,
37,
37,
37,
37,
37,
38,
38,
38,
38,
38,
38,
38,
39,
39,
39,
39,
39,
39,
39,
39,
39,
39,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
40,
41,
41,
41,
41,
41,
41,
41,
42,
42,
42,
42,
42,
42,
42,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
43,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
44,
45,
45,
45,
45,
45,
45,
45,
45,
45,
45,
45,
45,
45,
45,
45,
45,
46,
46,
46,
46,
46,
46,
46,
46,
46,
46,
46,
46,
46,
46,
47,
47,
47,
47,
47,
47,
47,
47,
47,
47,
47,
47,
47,
47,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
48,
49,
49,
49,
49,
49,
49,
49,
49,
49,
49,
49,
49,
49,
49,
49,
49,
50,
50,
50,
50,
50,
50,
50,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
51,
52,
52,
52,
52,
52,
52,
52,
52,
52,
52,
52,
52,
52,
52,
52,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
53,
54,
54,
54,
54,
54,
54,
54,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
55,
56,
56,
56,
56,
56,
56,
56,
56,
56,
56,
56,
56,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
57,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
58,
59,
59,
59,
59,
59,
59,
59,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
60,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
61,
62,
62,
62,
62,
62,
62,
62,
62,
62,
62,
62,
62,
62,
62,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
63,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
64,
65,
65,
65,
65,
65,
65,
65,
66,
66,
66,
66,
66,
66,
66,
66,
66,
66,
66,
67,
67,
67,
67,
67,
67,
67,
67,
67,
67,
67,
67,
67,
67,
67,
67,
68,
68,
68,
68,
68,
68,
68,
68,
68,
68,
68,
68,
68,
68,
68,
69,
69,
69,
69,
69,
69,
69,
69,
69,
69,
69,
69,
69,
69,
70,
70,
70,
70,
70,
70,
70,
71,
71,
71,
71,
71,
71,
71,
71,
71,
71,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
72,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
73,
74,
74,
74,
74,
74,
74,
74,
74,
74,
74,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
75,
76,
76,
76,
76,
76,
76,
76,
77,
77,
77,
77,
77,
77,
77,
77,
77,
77,
77,
77,
77,
77,
77,
77,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
78,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
79,
80,
80,
80,
80,
80,
80,
80,
80,
80,
80,
80,
80,
80,
80,
81,
81,
81,
81,
81,
81,
81,
81,
81,
81,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
82,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
83,
84,
84,
84,
84,
84,
84,
84,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
85,
86,
86,
86,
86,
86,
86,
86,
86,
86,
86,
86,
86,
86,
86,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
87,
88,
88,
88,
88,
88,
88,
88,
88,
88,
88,
88,
88,
88,
88,
89,
89,
89,
89,
89,
89,
89,
89,
89,
89,
89,
89,
90,
90,
90,
90,
90,
90,
90,
90,
90,
90,
90,
90,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
91,
92,
92,
92,
92,
92,
92,
92,
92,
92,
92,
92,
92,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
93,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
94,
95,
95,
95,
95,
95,
95,
95,
95,
95,
95,
95,
95,
95,
95,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
96,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
97,
98,
98,
98,
98,
98,
98,
98,
99,
99,
99,
99,
99,
99,
99,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
100,
101,
101,
101,
101,
101,
101,
101,
101,
101,
101,
101,
101,
101,
101,
101,
101,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
102,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
103,
104,
104,
104,
104,
104,
104,
104,
104,
104,
104,
105,
105,
105,
105,
105,
105,
105,
105,
105,
105,
105,
105,
106,
106,
106,
106,
106,
106,
106,
106,
106,
106,
106,
106,
106,
106,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
107,
108,
108,
108,
108,
108,
108,
108,
108,
108,
108,
108,
109,
109,
109,
109,
109,
109,
109,
109,
109,
109,
109,
109,
109,
109,
110,
110,
110,
110,
110,
110,
110,
110,
110,
110,
110,
110,
110,
110,
110,
110,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
111,
112,
112,
112,
112,
112,
112,
112,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
113,
114,
114,
114,
114,
114,
114,
114,
114,
114,
114,
114,
114,
114,
114,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
115,
116,
116,
116,
116,
116,
116,
116,
116,
116,
116,
116,
116,
117,
117,
117,
117,
117,
117,
117,
117,
117,
117,
117,
117,
117,
117,
118,
118,
118,
118,
118,
118,
118,
119,
119,
119,
119,
119,
119,
119,
119,
119,
119,
119,
119,
119,
119,
119,
119,
120,
120,
120,
120,
120,
120,
120,
120,
120,
120,
120,
121,
121,
121,
121,
121,
121,
121,
121,
121,
121,
121,
121,
121,
121,
122,
122,
122,
122,
122,
122,
122,
122,
122,
122,
122,
122,
122,
122,
122,
122,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
123,
124,
124,
124,
124,
124,
124,
124,
124,
124,
124,
125,
125,
125,
125,
125,
125,
125,
126,
126,
126,
126,
126,
126,
126,
127,
127,
127,
127,
127,
127,
127,
127,
127,
127,
127,
127,
127,
127,
127,
127,
128,
128,
128,
128,
128,
128,
128,
128,
128,
128,
128,
128,
128,
128,
128,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
129,
130,
130,
130,
130,
130,
130,
130,
130,
130,
130,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
131,
132,
132,
132,
132,
132,
132,
132,
132,
132,
132,
132,
132,
132,
132,
133,
133,
133,
133,
133,
133,
133,
133,
133,
133,
133,
133,
133,
133,
134,
134,
134,
134,
134,
134,
134,
134,
134,
134,
134,
134,
134,
134,
134,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
135,
136,
136,
136,
136,
136,
136,
136,
136,
136,
136,
137,
137,
137,
137,
137,
137,
137,
137,
137,
137,
137,
137,
137,
137,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
138,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
139,
140,
140,
140,
140,
140,
140,
140,
140,
140,
140,
140,
140,
140,
140,
140,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
141,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
142,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
143,
144,
144,
144,
144,
144,
144,
144,
144,
144,
144,
144,
144,
144,
144,
145,
145,
145,
145,
145,
145,
145,
145,
145,
145,
145,
145,
145,
145,
146,
146,
146,
146,
146,
146,
146,
146,
146,
146,
146,
146,
146,
146,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
147,
148,
148,
148,
148,
148,
148,
148,
149,
149,
149,
149,
149,
149,
149,
149,
149,
149,
149,
149,
150,
150,
150,
150,
150,
150,
150,
150,
150,
150,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
151,
152,
152,
152,
152,
152,
152,
152,
152,
152,
152,
152,
152,
152,
152,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
153,
154,
154,
154,
154,
154,
154,
154,
155,
155,
155,
155,
155,
155,
155,
155,
155,
155,
155,
155,
155,
155,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
156,
157,
157,
157,
157,
157,
157,
157,
157,
157,
157,
157,
157,
157,
157,
158,
158,
158,
158,
158,
158,
158,
158,
158,
158,
158,
158,
159,
159,
159,
159,
159,
159,
159,
159,
159,
159,
159,
159,
159,
159,
160,
160,
160,
160,
160,
160,
160,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
161,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
162,
163,
163,
163,
163,
163,
163,
163,
163,
163,
163,
163,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
164,
165,
165,
165,
165,
165,
165,
165,
166,
166,
166,
166,
166,
166,
166,
166,
166,
166,
166,
166,
166,
166,
166,
166,
167,
167,
167,
167,
167,
167,
167,
167,
167,
167,
167,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
168,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
169,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
170,
171,
171,
171,
171,
171,
171,
171;
	chainnames = 
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A",
"A";
	dynamicstate = 
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1,
1;
	nbspringsperparticle = 
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0;
}
